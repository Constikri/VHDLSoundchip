----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Wed Aug 18 14:23:38 2021
-- Parameters for CoreTimer
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant HDL_license : string( 1 to 1 ) := "O";
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 32;
end coreparameters;
