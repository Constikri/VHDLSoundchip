--------------------------------------------------------------------------------
-- Company: <Name>
--
-- File: dsp.vhd
-- File history:
--      <Revision number>: <Date>: <Comments>
--      <Revision number>: <Date>: <Comments>
--      <Revision number>: <Date>: <Comments>
--
-- Description: 
--
-- <Description here>
--
-- Targeted device: <Family::SmartFusion2> <Die::M2S010> <Package::256 VF>
-- Author: <Name>
--
--------------------------------------------------------------------------------

library IEEE;

use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

entity soundchip_hdl is
port (
    --<port_name> : <direction> <type>;
    --IN SPI
    -- OUT:
    OUT_0 : OUT std_logic;
    OUT_1 : OUT std_logic;
    OUT_2 : OUT std_logic;
    OUT_3 : OUT std_logic;
    OUT_4 : OUT std_logic;
    OUT_5 : OUT std_logic;
    OUT_6 : OUT std_logic;
    OUT_7 : OUT std_logic;
    OUT_8 : OUT std_logic;
    OUT_9 : OUT std_logic;
    OUT_10 : OUT std_logic;
    OUT_11 : OUT std_logic;
    OUT_12 : OUT std_logic;
    OUT_13 : OUT std_logic;
    OUT_14 : OUT std_logic;
    OUT_15 : OUT std_logic
);
end soundchip_hdl;
architecture architecture_soundchip_hdl of soundchip_hdl is
   -- signal, component etc. declarations

begin

   -- architecture body
end architecture_soundchip_hdl;
