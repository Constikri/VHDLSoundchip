----------------------------------------------------------------------
-- Created by SmartDesign Thu Aug 19 11:59:18 2021
-- Version: v2021.1 2021.1.0.17
----------------------------------------------------------------------

----------------------------------------------------------------------
-- Component Description (Tcl) 
----------------------------------------------------------------------
--# Exporting Component Description of CoreGPIO_C0 to TCL
--# Family: SmartFusion2
--# Part Number: M2S010-VF256
--# Create and Configure the core component CoreGPIO_C0
--create_and_configure_core -core_vlnv {Actel:DirectCore:CoreGPIO:3.0.120} -component_name {CoreGPIO_C0} -params {\
--"APB_WIDTH:32"  \
--"FIXED_CONFIG_0:false"  \
--"FIXED_CONFIG_1:false"  \
--"FIXED_CONFIG_2:false"  \
--"FIXED_CONFIG_3:false"  \
--"FIXED_CONFIG_4:false"  \
--"FIXED_CONFIG_5:false"  \
--"FIXED_CONFIG_6:false"  \
--"FIXED_CONFIG_7:false"  \
--"FIXED_CONFIG_8:false"  \
--"FIXED_CONFIG_9:false"  \
--"FIXED_CONFIG_10:false"  \
--"FIXED_CONFIG_11:false"  \
--"FIXED_CONFIG_12:false"  \
--"FIXED_CONFIG_13:false"  \
--"FIXED_CONFIG_14:false"  \
--"FIXED_CONFIG_15:false"  \
--"FIXED_CONFIG_16:false"  \
--"FIXED_CONFIG_17:false"  \
--"FIXED_CONFIG_18:false"  \
--"FIXED_CONFIG_19:false"  \
--"FIXED_CONFIG_20:false"  \
--"FIXED_CONFIG_21:false"  \
--"FIXED_CONFIG_22:false"  \
--"FIXED_CONFIG_23:false"  \
--"FIXED_CONFIG_24:false"  \
--"FIXED_CONFIG_25:false"  \
--"FIXED_CONFIG_26:false"  \
--"FIXED_CONFIG_27:false"  \
--"FIXED_CONFIG_28:false"  \
--"FIXED_CONFIG_29:false"  \
--"FIXED_CONFIG_30:false"  \
--"FIXED_CONFIG_31:false"  \
--"INT_BUS:0"  \
--"IO_INT_TYPE_0:7"  \
--"IO_INT_TYPE_1:7"  \
--"IO_INT_TYPE_2:7"  \
--"IO_INT_TYPE_3:7"  \
--"IO_INT_TYPE_4:7"  \
--"IO_INT_TYPE_5:7"  \
--"IO_INT_TYPE_6:7"  \
--"IO_INT_TYPE_7:7"  \
--"IO_INT_TYPE_8:7"  \
--"IO_INT_TYPE_9:7"  \
--"IO_INT_TYPE_10:7"  \
--"IO_INT_TYPE_11:7"  \
--"IO_INT_TYPE_12:7"  \
--"IO_INT_TYPE_13:7"  \
--"IO_INT_TYPE_14:7"  \
--"IO_INT_TYPE_15:7"  \
--"IO_INT_TYPE_16:7"  \
--"IO_INT_TYPE_17:7"  \
--"IO_INT_TYPE_18:7"  \
--"IO_INT_TYPE_19:7"  \
--"IO_INT_TYPE_20:7"  \
--"IO_INT_TYPE_21:7"  \
--"IO_INT_TYPE_22:7"  \
--"IO_INT_TYPE_23:7"  \
--"IO_INT_TYPE_24:7"  \
--"IO_INT_TYPE_25:7"  \
--"IO_INT_TYPE_26:7"  \
--"IO_INT_TYPE_27:7"  \
--"IO_INT_TYPE_28:7"  \
--"IO_INT_TYPE_29:7"  \
--"IO_INT_TYPE_30:7"  \
--"IO_INT_TYPE_31:7"  \
--"IO_NUM:32"  \
--"IO_TYPE_0:0"  \
--"IO_TYPE_1:0"  \
--"IO_TYPE_2:0"  \
--"IO_TYPE_3:0"  \
--"IO_TYPE_4:0"  \
--"IO_TYPE_5:0"  \
--"IO_TYPE_6:0"  \
--"IO_TYPE_7:0"  \
--"IO_TYPE_8:0"  \
--"IO_TYPE_9:0"  \
--"IO_TYPE_10:0"  \
--"IO_TYPE_11:0"  \
--"IO_TYPE_12:0"  \
--"IO_TYPE_13:0"  \
--"IO_TYPE_14:0"  \
--"IO_TYPE_15:0"  \
--"IO_TYPE_16:0"  \
--"IO_TYPE_17:0"  \
--"IO_TYPE_18:0"  \
--"IO_TYPE_19:0"  \
--"IO_TYPE_20:0"  \
--"IO_TYPE_21:0"  \
--"IO_TYPE_22:0"  \
--"IO_TYPE_23:0"  \
--"IO_TYPE_24:0"  \
--"IO_TYPE_25:0"  \
--"IO_TYPE_26:0"  \
--"IO_TYPE_27:0"  \
--"IO_TYPE_28:0"  \
--"IO_TYPE_29:0"  \
--"IO_TYPE_30:0"  \
--"IO_TYPE_31:0"  \
--"IO_VAL_0:0"  \
--"IO_VAL_1:0"  \
--"IO_VAL_2:0"  \
--"IO_VAL_3:0"  \
--"IO_VAL_4:0"  \
--"IO_VAL_5:0"  \
--"IO_VAL_6:0"  \
--"IO_VAL_7:0"  \
--"IO_VAL_8:0"  \
--"IO_VAL_9:0"  \
--"IO_VAL_10:0"  \
--"IO_VAL_11:0"  \
--"IO_VAL_12:0"  \
--"IO_VAL_13:0"  \
--"IO_VAL_14:0"  \
--"IO_VAL_15:0"  \
--"IO_VAL_16:0"  \
--"IO_VAL_17:0"  \
--"IO_VAL_18:0"  \
--"IO_VAL_19:0"  \
--"IO_VAL_20:0"  \
--"IO_VAL_21:0"  \
--"IO_VAL_22:0"  \
--"IO_VAL_23:0"  \
--"IO_VAL_24:0"  \
--"IO_VAL_25:0"  \
--"IO_VAL_26:0"  \
--"IO_VAL_27:0"  \
--"IO_VAL_28:0"  \
--"IO_VAL_29:0"  \
--"IO_VAL_30:0"  \
--"IO_VAL_31:0"  \
--"OE_TYPE:0"   }
--# Exporting Component Description of CoreGPIO_C0 to TCL done

----------------------------------------------------------------------
-- Libraries
----------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library smartfusion2;
use smartfusion2.all;
library COREGPIO_LIB;
use COREGPIO_LIB.all;
use COREGPIO_LIB.components.all;
----------------------------------------------------------------------
-- CoreGPIO_C0 entity declaration
----------------------------------------------------------------------
entity CoreGPIO_C0 is
    -- Port list
    port(
        -- Inputs
        GPIO_IN  : in  std_logic_vector(31 downto 0);
        PADDR    : in  std_logic_vector(7 downto 0);
        PCLK     : in  std_logic;
        PENABLE  : in  std_logic;
        PRESETN  : in  std_logic;
        PSEL     : in  std_logic;
        PWDATA   : in  std_logic_vector(31 downto 0);
        PWRITE   : in  std_logic;
        -- Outputs
        GPIO_OE  : out std_logic_vector(31 downto 0);
        GPIO_OUT : out std_logic_vector(31 downto 0);
        INT      : out std_logic_vector(31 downto 0);
        PRDATA   : out std_logic_vector(31 downto 0);
        PREADY   : out std_logic;
        PSLVERR  : out std_logic
        );
end CoreGPIO_C0;
----------------------------------------------------------------------
-- CoreGPIO_C0 architecture body
----------------------------------------------------------------------
architecture RTL of CoreGPIO_C0 is
----------------------------------------------------------------------
-- Component declarations
----------------------------------------------------------------------
-- CoreGPIO   -   Actel:DirectCore:CoreGPIO:3.0.120
-- using entity instantiation for component CoreGPIO
----------------------------------------------------------------------
-- Signal declarations
----------------------------------------------------------------------
signal APB_bif_PRDATA        : std_logic_vector(31 downto 0);
signal APB_bif_PREADY        : std_logic;
signal APB_bif_PSLVERR       : std_logic;
signal GPIO_OE_net_0         : std_logic_vector(31 downto 0);
signal GPIO_OUT_net_0        : std_logic_vector(31 downto 0);
signal INT_net_0             : std_logic_vector(31 downto 0);
signal INT_net_1             : std_logic_vector(31 downto 0);
signal GPIO_OUT_net_1        : std_logic_vector(31 downto 0);
signal GPIO_OE_net_1         : std_logic_vector(31 downto 0);
signal APB_bif_PRDATA_net_0  : std_logic_vector(31 downto 0);
signal APB_bif_PREADY_net_0  : std_logic;
signal APB_bif_PSLVERR_net_0 : std_logic;

begin
----------------------------------------------------------------------
-- Top level output port assignments
----------------------------------------------------------------------
 INT_net_1             <= INT_net_0;
 INT(31 downto 0)      <= INT_net_1;
 GPIO_OUT_net_1        <= GPIO_OUT_net_0;
 GPIO_OUT(31 downto 0) <= GPIO_OUT_net_1;
 GPIO_OE_net_1         <= GPIO_OE_net_0;
 GPIO_OE(31 downto 0)  <= GPIO_OE_net_1;
 APB_bif_PRDATA_net_0  <= APB_bif_PRDATA;
 PRDATA(31 downto 0)   <= APB_bif_PRDATA_net_0;
 APB_bif_PREADY_net_0  <= APB_bif_PREADY;
 PREADY                <= APB_bif_PREADY_net_0;
 APB_bif_PSLVERR_net_0 <= APB_bif_PSLVERR;
 PSLVERR               <= APB_bif_PSLVERR_net_0;
----------------------------------------------------------------------
-- Component instances
----------------------------------------------------------------------
-- CoreGPIO_C0_0   -   Actel:DirectCore:CoreGPIO:3.0.120
CoreGPIO_C0_0 : entity COREGPIO_LIB.CoreGPIO
    generic map( 
        APB_WIDTH       => ( 32 ),
        FAMILY          => ( 11 ),
        FIXED_CONFIG_0  => ( 0 ),
        FIXED_CONFIG_1  => ( 0 ),
        FIXED_CONFIG_2  => ( 0 ),
        FIXED_CONFIG_3  => ( 0 ),
        FIXED_CONFIG_4  => ( 0 ),
        FIXED_CONFIG_5  => ( 0 ),
        FIXED_CONFIG_6  => ( 0 ),
        FIXED_CONFIG_7  => ( 0 ),
        FIXED_CONFIG_8  => ( 0 ),
        FIXED_CONFIG_9  => ( 0 ),
        FIXED_CONFIG_10 => ( 0 ),
        FIXED_CONFIG_11 => ( 0 ),
        FIXED_CONFIG_12 => ( 0 ),
        FIXED_CONFIG_13 => ( 0 ),
        FIXED_CONFIG_14 => ( 0 ),
        FIXED_CONFIG_15 => ( 0 ),
        FIXED_CONFIG_16 => ( 0 ),
        FIXED_CONFIG_17 => ( 0 ),
        FIXED_CONFIG_18 => ( 0 ),
        FIXED_CONFIG_19 => ( 0 ),
        FIXED_CONFIG_20 => ( 0 ),
        FIXED_CONFIG_21 => ( 0 ),
        FIXED_CONFIG_22 => ( 0 ),
        FIXED_CONFIG_23 => ( 0 ),
        FIXED_CONFIG_24 => ( 0 ),
        FIXED_CONFIG_25 => ( 0 ),
        FIXED_CONFIG_26 => ( 0 ),
        FIXED_CONFIG_27 => ( 0 ),
        FIXED_CONFIG_28 => ( 0 ),
        FIXED_CONFIG_29 => ( 0 ),
        FIXED_CONFIG_30 => ( 0 ),
        FIXED_CONFIG_31 => ( 0 ),
        INT_BUS         => ( 0 ),
        IO_INT_TYPE_0   => ( 7 ),
        IO_INT_TYPE_1   => ( 7 ),
        IO_INT_TYPE_2   => ( 7 ),
        IO_INT_TYPE_3   => ( 7 ),
        IO_INT_TYPE_4   => ( 7 ),
        IO_INT_TYPE_5   => ( 7 ),
        IO_INT_TYPE_6   => ( 7 ),
        IO_INT_TYPE_7   => ( 7 ),
        IO_INT_TYPE_8   => ( 7 ),
        IO_INT_TYPE_9   => ( 7 ),
        IO_INT_TYPE_10  => ( 7 ),
        IO_INT_TYPE_11  => ( 7 ),
        IO_INT_TYPE_12  => ( 7 ),
        IO_INT_TYPE_13  => ( 7 ),
        IO_INT_TYPE_14  => ( 7 ),
        IO_INT_TYPE_15  => ( 7 ),
        IO_INT_TYPE_16  => ( 7 ),
        IO_INT_TYPE_17  => ( 7 ),
        IO_INT_TYPE_18  => ( 7 ),
        IO_INT_TYPE_19  => ( 7 ),
        IO_INT_TYPE_20  => ( 7 ),
        IO_INT_TYPE_21  => ( 7 ),
        IO_INT_TYPE_22  => ( 7 ),
        IO_INT_TYPE_23  => ( 7 ),
        IO_INT_TYPE_24  => ( 7 ),
        IO_INT_TYPE_25  => ( 7 ),
        IO_INT_TYPE_26  => ( 7 ),
        IO_INT_TYPE_27  => ( 7 ),
        IO_INT_TYPE_28  => ( 7 ),
        IO_INT_TYPE_29  => ( 7 ),
        IO_INT_TYPE_30  => ( 7 ),
        IO_INT_TYPE_31  => ( 7 ),
        IO_NUM          => ( 32 ),
        IO_TYPE_0       => ( 0 ),
        IO_TYPE_1       => ( 0 ),
        IO_TYPE_2       => ( 0 ),
        IO_TYPE_3       => ( 0 ),
        IO_TYPE_4       => ( 0 ),
        IO_TYPE_5       => ( 0 ),
        IO_TYPE_6       => ( 0 ),
        IO_TYPE_7       => ( 0 ),
        IO_TYPE_8       => ( 0 ),
        IO_TYPE_9       => ( 0 ),
        IO_TYPE_10      => ( 0 ),
        IO_TYPE_11      => ( 0 ),
        IO_TYPE_12      => ( 0 ),
        IO_TYPE_13      => ( 0 ),
        IO_TYPE_14      => ( 0 ),
        IO_TYPE_15      => ( 0 ),
        IO_TYPE_16      => ( 0 ),
        IO_TYPE_17      => ( 0 ),
        IO_TYPE_18      => ( 0 ),
        IO_TYPE_19      => ( 0 ),
        IO_TYPE_20      => ( 0 ),
        IO_TYPE_21      => ( 0 ),
        IO_TYPE_22      => ( 0 ),
        IO_TYPE_23      => ( 0 ),
        IO_TYPE_24      => ( 0 ),
        IO_TYPE_25      => ( 0 ),
        IO_TYPE_26      => ( 0 ),
        IO_TYPE_27      => ( 0 ),
        IO_TYPE_28      => ( 0 ),
        IO_TYPE_29      => ( 0 ),
        IO_TYPE_30      => ( 0 ),
        IO_TYPE_31      => ( 0 ),
        IO_VAL_0        => ( 0 ),
        IO_VAL_1        => ( 0 ),
        IO_VAL_2        => ( 0 ),
        IO_VAL_3        => ( 0 ),
        IO_VAL_4        => ( 0 ),
        IO_VAL_5        => ( 0 ),
        IO_VAL_6        => ( 0 ),
        IO_VAL_7        => ( 0 ),
        IO_VAL_8        => ( 0 ),
        IO_VAL_9        => ( 0 ),
        IO_VAL_10       => ( 0 ),
        IO_VAL_11       => ( 0 ),
        IO_VAL_12       => ( 0 ),
        IO_VAL_13       => ( 0 ),
        IO_VAL_14       => ( 0 ),
        IO_VAL_15       => ( 0 ),
        IO_VAL_16       => ( 0 ),
        IO_VAL_17       => ( 0 ),
        IO_VAL_18       => ( 0 ),
        IO_VAL_19       => ( 0 ),
        IO_VAL_20       => ( 0 ),
        IO_VAL_21       => ( 0 ),
        IO_VAL_22       => ( 0 ),
        IO_VAL_23       => ( 0 ),
        IO_VAL_24       => ( 0 ),
        IO_VAL_25       => ( 0 ),
        IO_VAL_26       => ( 0 ),
        IO_VAL_27       => ( 0 ),
        IO_VAL_28       => ( 0 ),
        IO_VAL_29       => ( 0 ),
        IO_VAL_30       => ( 0 ),
        IO_VAL_31       => ( 0 ),
        OE_TYPE         => ( 0 )
        )
    port map( 
        -- Inputs
        PRESETN  => PRESETN,
        PCLK     => PCLK,
        PSEL     => PSEL,
        PENABLE  => PENABLE,
        PWRITE   => PWRITE,
        PADDR    => PADDR,
        PWDATA   => PWDATA,
        GPIO_IN  => GPIO_IN,
        -- Outputs
        PSLVERR  => APB_bif_PSLVERR,
        PREADY   => APB_bif_PREADY,
        PRDATA   => APB_bif_PRDATA,
        INT      => INT_net_0,
        INT_OR   => OPEN,
        GPIO_OUT => GPIO_OUT_net_0,
        GPIO_OE  => GPIO_OE_net_0 
        );

end RTL;
