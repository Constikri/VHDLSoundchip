--  Copyright 2011 Actel Corporation.  All rights reserved.
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
-- ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
-- Revision Information:
-- SVN Revision Information:
-- SVN $Revision: 4805 $
library ieEE;
use IEee.STD_lOGIc_1164.all;
use IeeE.stD_logIC_ariTH.all;
use ieeE.STd_lOGic_UNSignED.all;
use ieeE.sTD_loGIC_mISC.all;
entity CHTOLSRAMoo1 is
generic (uSRam_NUM_lOCAtioNS_dwIDth32: iNTEger := 128); port (CHTOLSRAMLO1: in STd_lOGIc_VECtor(7 downto 0);
CHTOLSRAMio1: out STd_lOGic_VECtoR(7 downto 0);
WEn: in sTD_logIC;
reN: in STD_loGIc;
CHTOLSRAMOL1: in sTD_loGIC_veCTor(15 downto 0);
CHTOLSRAMLl1: in Std_LOgic_VectOR(15 downto 0);
clK: in Std_LOgic;
CHTOLSRAMIL1: in STd_lOGIc;
CHTOLSRAMoi1: out sTD_loGIC);
end entity CHTOLSRAMOO1;

architecture CHTOLSRAMO of CHTOLSRAMOO1 is

component RAM64x18
port (a_Dout: out STd_LOGic_VEctoR(17 downto 0);
B_doUT: out sTD_logIC_veCTOr(17 downto 0);
A_adDr_cLk: in std_LoGiC;
b_Addr_CLk: in STD_lOGIc;
A_addR_en: in sTD_loGIC;
B_AddR_En: in stD_LogiC;
a_aDDR_lAT: in STD_loGIC;
B_Addr_Lat: in stD_logIC;
A_adDR_arST_n: in STD_loGIC;
B_addR_Arst_N: in Std_LOgic;
a_ADDr_sRSt_n: in std_LogiC;
B_AddR_Srst_N: in std_LOgiC;
a_DoUT_clK: in std_LOgiC;
b_Dout_CLk: in stD_LogIC;
a_DOut_EN: in std_LOgiC;
b_Dout_EN: in std_LOgic;
a_DOut_LAt: in stD_logIC;
b_DOUt_LAT: in std_LOgic;
A_douT_Arst_N: in stD_LogIC;
b_DOut_ARst_N: in STd_lOGIc;
A_douT_SrsT_N: in stD_LogIC;
b_DOut_SRSt_n: in stD_LogiC;
A_addR: in Std_LOgic_VEctOR(9 downto 0);
b_ADdr: in stD_LogiC_vecTOR(9 downto 0);
a_WIDth: in stD_LogiC_vecTOR(2 downto 0);
B_WidTH: in stD_logIC_vecTOr(2 downto 0);
A_blk: in STd_lOGic_VECtor(1 downto 0);
B_blK: in Std_LOGic_VEctoR(1 downto 0);
a_EN: in Std_LOGic;
b_EN: in sTD_loGIC;
C_clK: in stD_LogiC;
c_bLK: in STD_lOGIc_vECTor(1 downto 0);
c_DIN: in std_LogiC_VecTOR(17 downto 0);
C_en: in stD_logIC;
C_adDR: in Std_LOGic_VEctoR(9 downto 0);
c_Wen: in Std_LOGic;
c_WIdth: in STd_lOGIc_vECtor(2 downto 0);
BUsy: out Std_LOGic;
Sii_LOCk: in sTD_loGIC);
end component;

signal CHTOLSRAMl1LL: std_LogiC_VecTOR(13 downto 6);

signal WidtH0: STD_lOGIc_vECTor(2 downto 0);

signal WIDth1: sTD_logIC_veCTOr(2 downto 0);

signal WidtH2: sTD_loGIC_veCTOr(2 downto 0);

signal CHTOLSRAMi1LL: STd_lOGic_VECtor(2 downto 0);

signal CHTOLSRAMOoil: sTD_logIC_veCTOr(2 downto 0);

signal CHTOLSRAMloiL: STd_lOGIc_vECtor(2 downto 0);

signal CHTOLSRAMiOIL: stD_logIC_vecTOr(2 downto 0);

signal CHTOLSRAMOliL: sTD_logIC_veCTOr(2 downto 0);

signal CHTOLSRAMlliL: STd_lOGIc_vECtor(2 downto 0);

signal CHTOLSRAMiLIL: Std_LOGic_VEctoR(2 downto 0);

signal CHTOLSRAMOIil: std_LOgiC_VectOR(2 downto 0);

signal CHTOLSRAMliIL: STD_lOGIc_vECtor(2 downto 0);

signal CHTOLSRAMiiiL: STd_LOGic_VECtoR(2 downto 0);

signal CHTOLSRAMO0il: sTD_loGIC_veCTor(2 downto 0);

signal CHTOLSRAMl0iL: STD_loGIC_vECTor(2 downto 0);

signal CHTOLSRAMi0IL: stD_LogiC_vecTOR(2 downto 0);

signal CHTOLSRAMO1il: sTD_loGIC_veCTOr(2 downto 0);

signal CHTOLSRAML1il: stD_logIC_vecTOr(2 downto 0);

signal CHTOLSRAMi1iL: Std_LOgic;

signal CHTOLSRAMoO0L: stD_LogiC;

signal CHTOLSRAMLo0l: STd_lOGIc;

signal CHTOLSRAMio0L: Std_LOgic;

signal CHTOLSRAMOL0l: sTD_loGIC;

signal CHTOLSRAMLl0l: STd_LOGic;

signal CHTOLSRAMil0L: std_LOgiC;

signal CHTOLSRAMoI0L: stD_LogIC;

signal CHTOLSRAMli0L: std_LogiC;

signal CHTOLSRAMII0l: STd_lOGIc;

signal CHTOLSRAMO00l: STd_lOGic;

signal CHTOLSRAMl00L: Std_LOGic;

signal CHTOLSRAMI00l: sTD_logIC;

signal CHTOLSRAMo10L: Std_LOgic;

signal CHTOLSRAMl10l: sTD_loGIC;

signal CHTOLSRAMI10L: Std_LOgic;

signal CHTOLSRAMOo1l: Std_LOGic;

signal CHTOLSRAMlO1L: stD_LOGIc;

signal CHTOLSRAMio1L: stD_LogiC;

signal CHTOLSRAMol1L: Std_LOGic;

signal CHTOLSRAMlL1L: sTD_loGIC;

signal CHTOLSRAMil1L: std_LOgiC;

signal CHTOLSRAMOI1l: STD_lOGIc;

signal CHTOLSRAMli1L: Std_LOgic;

signal CHTOLSRAMII1l: STD_loGIC;

signal CHTOLSRAMo01L: STd_LOGic;

signal CHTOLSRAMl01L: std_LOgic;

signal CHTOLSRAMI01l: sTD_logIC;

signal CHTOLSRAMo11L: Std_LOgic;

signal CHTOLSRAML11l: sTD_loGIC;

signal CHTOLSRAMi11L: Std_LOGic;

signal CHTOLSRAMOOoi: sTD_loGIC;

signal CHTOLSRAMloOI: stD_LogiC;

signal CHTOLSRAMIOoi: sTD_logIC;

signal CHTOLSRAMolOI: Std_LOGic;

signal CHTOLSRAMlLOi: std_LogiC;

signal CHTOLSRAMilOI: STD_lOGIc_vECTor(17 downto 0);

signal CHTOLSRAMoiOI: Std_LOgic_VEctoR(17 downto 0);

signal CHTOLSRAMLIoi: std_LOgiC_VectOR(17 downto 0);

signal CHTOLSRAMIioI: Std_LOgic_VectOR(17 downto 0);

signal CHTOLSRAMo0oI: sTD_loGIC_veCTor(17 downto 0);

signal CHTOLSRAMl0OI: STD_loGIc_vECTor(17 downto 0);

signal CHTOLSRAMi0OI: STD_loGIc_vECTor(17 downto 0);

signal CHTOLSRAMO1Oi: sTD_loGIC_veCTOr(17 downto 0);

signal CHTOLSRAML1Oi: std_LogiC_VecTOR(17 downto 0);

signal CHTOLSRAMI1Oi: std_LOgiC_VectOR(17 downto 0);

signal CHTOLSRAMOoli: stD_LogiC_vecTOR(17 downto 0);

signal CHTOLSRAMLolI: sTD_loGIC_veCTor(17 downto 0);

signal CHTOLSRAMIOli: std_LogiC_VecTOR(17 downto 0);

signal CHTOLSRAMOLli: std_LogiC_VecTOR(17 downto 0);

signal CHTOLSRAMLLli: std_LOgic_VectOR(17 downto 0);

signal CHTOLSRAMILli: std_LogiC_VectOR(17 downto 0);

signal CHTOLSRAMoiLI: STd_lOGIc_vECtor(17 downto 0);

signal CHTOLSRAMLili: sTD_loGIC_veCTOr(17 downto 0);

signal CHTOLSRAMIIli: Std_LOgic_VEctoR(17 downto 0);

signal CHTOLSRAMO0li: stD_LogIC_vecTOR(17 downto 0);

signal CHTOLSRAML0li: stD_logIC_vecTOr(17 downto 0);

signal CHTOLSRAMI0Li: Std_LOGic_VEctoR(17 downto 0);

signal CHTOLSRAMo1LI: STD_lOGIc_vECTor(17 downto 0);

signal CHTOLSRAML1Li: std_LOgiC_VectOR(17 downto 0);

signal CHTOLSRAMi1lI: stD_LogIC_vecTOr(17 downto 0);

signal CHTOLSRAMOOIi: Std_LOgic_VectOR(17 downto 0);

signal CHTOLSRAMLoii: sTD_logIC_veCTOr(17 downto 0);

signal CHTOLSRAMioiI: Std_LOgic_VEctoR(17 downto 0);

signal CHTOLSRAMoliI: sTD_loGIC_veCTOr(17 downto 0);

signal CHTOLSRAMLlii: stD_logIC_veCTOr(17 downto 0);

signal CHTOLSRAMilII: STD_loGIC_vECTor(17 downto 0);

signal CHTOLSRAMOiii: stD_logIC_vecTOr(17 downto 0);

signal CHTOLSRAMLIii: std_LogiC_VecTOR(17 downto 0);

signal CHTOLSRAMIIii: stD_logIC_vecTOr(17 downto 0);

signal CHTOLSRAMo0Ii: Std_LOgic_VectOR(17 downto 0);

signal CHTOLSRAML0ii: std_LogiC_VecTOR(17 downto 0);

signal CHTOLSRAMI0ii: stD_logIC_vecTOr(9 downto 0);

signal CHTOLSRAMO1ii: std_LogiC_VecTOR(9 downto 0);

signal CHTOLSRAML1ii: stD_LogiC_vecTOR(9 downto 0);

signal CHTOLSRAMi1iI: sTD_loGIC_veCTor(9 downto 0);

signal CHTOLSRAMOo0i: sTD_logIC_veCTOr(9 downto 0);

signal CHTOLSRAMLo0I: sTD_logIC_veCTOr(9 downto 0);

signal CHTOLSRAMiO0I: Std_LOGic_VEctOR(9 downto 0);

signal CHTOLSRAMOL0i: Std_LOgic_VectOR(9 downto 0);

signal CHTOLSRAMlL0i: stD_LogiC_vecTOR(9 downto 0);

signal CHTOLSRAMil0I: STd_lOGic_VECtor(9 downto 0);

signal CHTOLSRAMoI0i: Std_LOGic_VEctoR(9 downto 0);

signal CHTOLSRAMLI0i: std_LOgiC_VectOR(9 downto 0);

signal CHTOLSRAMII0i: stD_LogIC_vecTOr(9 downto 0);

signal CHTOLSRAMO00i: stD_LogIC_vecTOr(9 downto 0);

signal CHTOLSRAML00I: stD_logIC_veCTOr(9 downto 0);

signal CHTOLSRAMi00I: STd_lOGIc_VECtor(9 downto 0);

signal CHTOLSRAMo10I: Std_LOGic_VEctoR(9 downto 0);

signal CHTOLSRAMl10I: STD_lOGIc_vECTor(9 downto 0);

signal CHTOLSRAMI10i: std_LogiC_VecTOR(9 downto 0);

signal CHTOLSRAMOO1i: Std_LOGic_VEctoR(9 downto 0);

signal CHTOLSRAMlO1I: STd_lOGIc_VECtor(9 downto 0);

signal CHTOLSRAMiO1I: STd_lOGIc_VECtor(9 downto 0);

signal CHTOLSRAMol1I: STd_lOGic_VECtoR(9 downto 0);

signal CHTOLSRAMLL1i: std_LogiC_VecTOR(9 downto 0);

signal CHTOLSRAMil1I: sTD_loGIC_veCTOr(9 downto 0);

signal CHTOLSRAMOi1i: stD_logIC_vecTOr(9 downto 0);

signal CHTOLSRAMLI1i: Std_LOgic_VectOR(9 downto 0);

signal CHTOLSRAMiI1I: STd_lOGIc_VECtor(9 downto 0);

signal CHTOLSRAMo01I: STd_lOGic_VECtor(9 downto 0);

signal CHTOLSRAMl01I: Std_LOgic_VectOR(9 downto 0);

signal CHTOLSRAMI01i: Std_LOgic_VectOR(9 downto 0);

signal CHTOLSRAMo11I: sTD_loGIC_veCTor(9 downto 0);

signal CHTOLSRAML11i: stD_LogiC_vecTOR(9 downto 0);

signal CHTOLSRAMi11I: STd_lOGic_VECtor(9 downto 0);

signal CHTOLSRAMooO0: STd_lOGic_VECtor(9 downto 0);

signal CHTOLSRAMlOO0: STd_LOGic_VECtoR(9 downto 0);

signal CHTOLSRAMI111: STd_LOGic_VECtoR(1 downto 0);

signal CHTOLSRAMOOOol: stD_LogIC_vecTOr(1 downto 0);

signal CHTOLSRAMLoooL: stD_logIC;

signal CHTOLSRAMioOOL: sTD_loGIC;

signal CHTOLSRAMoloOL: stD_LogIC;

signal CHTOLSRAMLLOol: STd_lOGIc;

signal CHTOLSRAMilOOl: STD_lOGIc;

signal CHTOLSRAMoioOL: stD_logIC;

signal CHTOLSRAMlioOL: Std_LOgic;

signal CHTOLSRAMIioOL: sTD_logIC;

signal CHTOLSRAMO0ool: Std_LOGic;

signal CHTOLSRAMl0OOL: sTD_loGIC;

signal CHTOLSRAMi0OOL: sTD_loGIC;

signal CHTOLSRAMO1Ool: STd_lOGIc;

signal CHTOLSRAMl1oOL: stD_logIC;

signal CHTOLSRAMI1ool: Std_LOgic;

signal CHTOLSRAMooLOl: STD_loGIC;

signal CHTOLSRAMLOlol: STd_lOGIc;

signal CHTOLSRAMIOlol: Std_LOGic;

signal CHTOLSRAMolLOL: stD_logIC;

signal CHTOLSRAMill0: STD_loGIc_vECTor(7 downto 0);

signal CHTOLSRAMLLlol: Std_LOgic;

begin
CHTOLSRAMIO1 <= CHTOLSRAMILl0;
CHTOLSRAMOi1 <= CHTOLSRAMLLloL;
process (CLk,CHTOLSRAMiL1)
begin
if (not CHTOLSRAMIL1 = '1') then
CHTOLSRAMl1LL(13 downto 6) <= "00000000";
elsif (Clk'evENT and clk = '1') then
CHTOLSRAML1lL(13 downto 6) <= CHTOLSRAMLL1(13 downto 6);
end if;
end process;
process (CHTOLSRAMLo1,CHTOLSRAMi1iL,CHTOLSRAMOo0l,CHTOLSRAMLO0l,CHTOLSRAMio0L,CHTOLSRAMOL0l,CHTOLSRAMll0L,CHTOLSRAML1ll,CHTOLSRAMll1,CHTOLSRAMOLii,CHTOLSRAMlLII,CHTOLSRAMilII,CHTOLSRAMOIii,CHTOLSRAMlIII,CHTOLSRAMIIii,wen,CHTOLSRAMo0iI,CHTOLSRAML0ii,CHTOLSRAMiiLI,CHTOLSRAMO0Li,CHTOLSRAMl0lI,CHTOLSRAMi0LI,CHTOLSRAMO1li,CHTOLSRAMl1LI,CHTOLSRAMI1Li,CHTOLSRAMoOIi,CHTOLSRAMLOii,CHTOLSRAMioII,CHTOLSRAMOL1)
variable CHTOLSRAMLIL0: std_LogiC_VectOR(2 downto 0);
variable CHTOLSRAMIIL0: STD_loGIC_veCTor(2 downto 0);
variable CHTOLSRAMO0l0: Std_LOgic_VectOR(2 downto 0);
variable CHTOLSRAMl0L0: Std_LOGic_VEctoR(2 downto 0);
variable CHTOLSRAMI0l0: Std_LOgic_VectOR(2 downto 0);
variable CHTOLSRAMo1L0: STd_lOGIc_vECtor(2 downto 0);
variable CHTOLSRAML1l0: STd_lOGic_VECtor(2 downto 0);
variable CHTOLSRAMi1L0: STd_lOGic_VECtor(2 downto 0);
variable CHTOLSRAMOOI0: Std_LOgic_VectOR(2 downto 0);
variable CHTOLSRAMLOi0: std_LOgiC_VectOR(2 downto 0);
variable CHTOLSRAMIOi0: std_LOgic_VectOR(2 downto 0);
variable CHTOLSRAMoli0: Std_LOgic_VectOR(2 downto 0);
variable CHTOLSRAMlLI0: STd_lOGic_VECtor(2 downto 0);
variable CHTOLSRAMiLI0: Std_LOGic_VEctoR(2 downto 0);
variable CHTOLSRAMoII0: STd_LOGic_VECtoR(2 downto 0);
variable CHTOLSRAMlII0: STd_lOGIc_vECtor(2 downto 0);
variable CHTOLSRAMiiI0: STD_loGIC_vECTor(2 downto 0);
variable CHTOLSRAMo0I0: STd_lOGIc_VECtor(2 downto 0);
variable CHTOLSRAMiLLOl: STd_lOGIc;
variable CHTOLSRAMOIloL: std_LOgic;
variable CHTOLSRAMlilOL: stD_LogIC;
variable CHTOLSRAMiILOl: STD_lOGIc;
variable CHTOLSRAMO0lol: STd_lOGic;
variable CHTOLSRAMl0lOL: stD_logIC;
variable CHTOLSRAMi0Lol: Std_LOGic;
variable CHTOLSRAMo1lOL: stD_logIC;
variable CHTOLSRAMl1lOL: STd_LOGic;
variable CHTOLSRAMi1lOL: sTD_logIC;
variable CHTOLSRAMOoioL: stD_LogiC;
variable CHTOLSRAMLOIol: STd_lOGIc;
variable CHTOLSRAMIOiol: Std_LOGic;
variable CHTOLSRAMolIOl: STD_loGIc;
variable CHTOLSRAMLLioL: std_LOgiC;
variable CHTOLSRAMilIOL: stD_logIC;
variable CHTOLSRAMOIIol: STd_lOGIc;
variable CHTOLSRAMliiOL: stD_LogIC;
variable CHTOLSRAMIIIol: STd_LOGic;
variable CHTOLSRAMo0IOL: sTD_loGIC;
variable CHTOLSRAML0ioL: Std_LOgic;
variable CHTOLSRAMi0iOL: stD_LogiC;
variable CHTOLSRAMo1IOl: STD_lOGIc;
variable CHTOLSRAML1ioL: std_LogiC;
variable CHTOLSRAMI1Iol: STD_lOGIc;
variable CHTOLSRAMoo0OL: stD_logIC;
variable CHTOLSRAMLO0ol: STd_lOGIc;
variable CHTOLSRAMio0Ol: sTD_loGIC;
variable CHTOLSRAMol0Ol: STD_loGIC;
variable CHTOLSRAMLl0oL: std_LOgiC;
variable CHTOLSRAMIL0ol: Std_LOGic;
variable CHTOLSRAMoi0OL: stD_logIC;
variable CHTOLSRAMlI0ol: STd_lOGIc;
variable CHTOLSRAMII0oL: Std_LOgic;
variable CHTOLSRAMo00OL: sTD_loGIC;
variable CHTOLSRAMl00ol: stD_LogiC_vecTOR(17 downto 0);
variable CHTOLSRAMi00OL: Std_LOGic_VEctoR(17 downto 0);
variable CHTOLSRAMO10ol: STd_lOGIc_VECtor(17 downto 0);
variable CHTOLSRAMl10Ol: stD_logIC_vecTOr(17 downto 0);
variable CHTOLSRAMi10Ol: std_LogiC_VecTOR(17 downto 0);
variable CHTOLSRAMoo1OL: STD_lOGIc_vECTor(17 downto 0);
variable CHTOLSRAMlO1ol: stD_logIC_vecTOr(17 downto 0);
variable CHTOLSRAMIO1oL: STD_loGIC_veCTor(17 downto 0);
variable CHTOLSRAMol1OL: Std_LOgic_VectOR(17 downto 0);
variable CHTOLSRAMLL1oL: sTD_loGIC_veCTOr(17 downto 0);
variable CHTOLSRAMIL1ol: stD_logIC_vecTOR(17 downto 0);
variable CHTOLSRAMoi1OL: std_LogiC_VectOR(17 downto 0);
variable CHTOLSRAMLi1oL: sTD_loGIC_veCTOr(17 downto 0);
variable CHTOLSRAMiI1Ol: std_LOgic_VectOR(17 downto 0);
variable CHTOLSRAMO01ol: sTD_logIC_veCTOr(17 downto 0);
variable CHTOLSRAML01oL: STD_loGIc_vECTor(17 downto 0);
variable CHTOLSRAMI01ol: sTD_logIC_veCTOr(17 downto 0);
variable CHTOLSRAMO11ol: sTD_logIC_veCTOr(17 downto 0);
variable CHTOLSRAMl11Ol: Std_LOgic_VEctoR(9 downto 0);
variable CHTOLSRAMI11ol: stD_LogIC_vecTOR(9 downto 0);
variable CHTOLSRAMoOOLl: std_LogiC_VecTOR(9 downto 0);
variable CHTOLSRAMloOLL: STd_lOGIc_VECtor(9 downto 0);
variable CHTOLSRAMIoolL: sTD_loGIC_veCTOr(9 downto 0);
variable CHTOLSRAMOlolL: STD_lOGIc_vECTor(9 downto 0);
variable CHTOLSRAMlLOLl: stD_LogiC_VecTOR(9 downto 0);
variable CHTOLSRAMIlolL: STD_lOGIc_vECTor(9 downto 0);
variable CHTOLSRAMoIOll: stD_LogiC_vecTOR(9 downto 0);
variable CHTOLSRAMlIOll: stD_LogiC_vecTOR(9 downto 0);
variable CHTOLSRAMIioLL: STd_lOGIc_vECtor(9 downto 0);
variable CHTOLSRAMO0olL: sTD_logIC_veCTOr(9 downto 0);
variable CHTOLSRAMl0OLL: stD_LogiC_vecTOR(9 downto 0);
variable CHTOLSRAMi0OLl: std_LogiC_VectOR(9 downto 0);
variable CHTOLSRAMO1oll: stD_LogIC_vecTOR(9 downto 0);
variable CHTOLSRAMl1OLl: std_LogiC_VectOR(9 downto 0);
variable CHTOLSRAMI1oll: sTD_loGIC_veCTOr(9 downto 0);
variable CHTOLSRAMooLLl: stD_LogiC_vecTOR(9 downto 0);
variable CHTOLSRAMloLLL: Std_LOGic_VEctor(9 downto 0);
variable CHTOLSRAMiOLLl: stD_logIC_vecTOR(9 downto 0);
variable CHTOLSRAMOllLL: Std_LOGic_VEctoR(9 downto 0);
variable CHTOLSRAMLlllL: STD_lOGIc_vECTor(9 downto 0);
variable CHTOLSRAMilLLL: Std_LOgic_VectOR(9 downto 0);
variable CHTOLSRAMOIlll: stD_logIC_vecTOR(9 downto 0);
variable CHTOLSRAMlILLl: sTD_loGIC_veCTOr(9 downto 0);
variable CHTOLSRAMiiLLL: Std_LOGic_VECtoR(9 downto 0);
variable CHTOLSRAMo0LLl: Std_LOgic_VEctoR(9 downto 0);
variable CHTOLSRAML0llL: STD_loGIC_vECTor(9 downto 0);
variable CHTOLSRAMi0lLL: Std_LOGic_VEctoR(9 downto 0);
variable CHTOLSRAMO1Lll: STD_loGIC_vECTor(9 downto 0);
variable CHTOLSRAMl1LLl: Std_LOgic_VEctoR(9 downto 0);
variable CHTOLSRAMI1lll: stD_logIC_vecTOR(9 downto 0);
variable CHTOLSRAMOoilL: STd_lOGIc_vECTor(9 downto 0);
variable CHTOLSRAMLoilL: STD_loGIC_veCTor(9 downto 0);
variable CHTOLSRAMioILl: Std_LOgic_VectOR(9 downto 0);
variable CHTOLSRAMOLill: stD_logIC_vecTOr(9 downto 0);
variable CHTOLSRAMlLILl: std_LOgic_VectOR(1 downto 0);
variable CHTOLSRAMILIll: stD_logIC_vecTOR(1 downto 0);
variable CHTOLSRAMOiilL: STD_lOGIc_vECTor(7 downto 0);
variable CHTOLSRAMlIIll: stD_LogiC_vecTOR(5 downto 0);
variable CHTOLSRAMIIilL: STd_lOGic_VECtor(2 downto 0);
begin
CHTOLSRAMLIl0 := "000";
CHTOLSRAMiiL0 := "000";
CHTOLSRAMO0l0 := "000";
CHTOLSRAML0l0 := "000";
CHTOLSRAMI0l0 := "000";
CHTOLSRAMo1L0 := "000";
CHTOLSRAMl1L0 := "000";
CHTOLSRAMI1l0 := "000";
CHTOLSRAMooi0 := "000";
CHTOLSRAMLOi0 := "000";
CHTOLSRAMIOi0 := "000";
CHTOLSRAMolI0 := "000";
CHTOLSRAMlli0 := "000";
CHTOLSRAMILi0 := "000";
CHTOLSRAMoii0 := "000";
CHTOLSRAMLIi0 := "000";
CHTOLSRAMiiI0 := "000";
CHTOLSRAMo0I0 := "000";
CHTOLSRAMILlol := '0';
CHTOLSRAMoILOl := '0';
CHTOLSRAMLiloL := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMO0Lol := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAMo1LOl := '0';
CHTOLSRAML1loL := '0';
CHTOLSRAMI1loL := '0';
CHTOLSRAMoOIol := '0';
CHTOLSRAMloiOL := '0';
CHTOLSRAMIoioL := '0';
CHTOLSRAMOlioL := '0';
CHTOLSRAMLLiol := '0';
CHTOLSRAMILiol := '0';
CHTOLSRAMOIIol := '0';
CHTOLSRAMLiioL := '0';
CHTOLSRAMIIioL := '0';
CHTOLSRAMO0iol := '0';
CHTOLSRAML0Iol := '0';
CHTOLSRAMI0iol := '0';
CHTOLSRAMO1Iol := '0';
CHTOLSRAMl1Iol := '0';
CHTOLSRAMi1IOl := '0';
CHTOLSRAMoO0Ol := '0';
CHTOLSRAMLo0OL := '0';
CHTOLSRAMIo0oL := '0';
CHTOLSRAMoL0ol := '0';
CHTOLSRAMll0OL := '0';
CHTOLSRAMIL0ol := '0';
CHTOLSRAMoI0ol := '0';
CHTOLSRAMLI0ol := '0';
CHTOLSRAMii0OL := '0';
CHTOLSRAMO00ol := '0';
CHTOLSRAML00ol := "000000000000000000";
CHTOLSRAMI00ol := "000000000000000000";
CHTOLSRAMo10Ol := "000000000000000000";
CHTOLSRAML10oL := "000000000000000000";
CHTOLSRAMI10oL := "000000000000000000";
CHTOLSRAMOo1oL := "000000000000000000";
CHTOLSRAMLo1oL := "000000000000000000";
CHTOLSRAMIO1ol := "000000000000000000";
CHTOLSRAMol1Ol := "000000000000000000";
CHTOLSRAMlL1Ol := "000000000000000000";
CHTOLSRAMiL1Ol := "000000000000000000";
CHTOLSRAMoI1Ol := "000000000000000000";
CHTOLSRAMli1OL := "000000000000000000";
CHTOLSRAMII1oL := "000000000000000000";
CHTOLSRAMo01ol := "000000000000000000";
CHTOLSRAML01ol := "000000000000000000";
CHTOLSRAMI01ol := "000000000000000000";
CHTOLSRAMO11ol := "000000000000000000";
CHTOLSRAMl11ol := "0000000000";
CHTOLSRAMI11oL := "0000000000";
CHTOLSRAMoOOLl := "0000000000";
CHTOLSRAMLOoll := "0000000000";
CHTOLSRAMioOLL := "0000000000";
CHTOLSRAMoLOLl := "0000000000";
CHTOLSRAMLLoll := "0000000000";
CHTOLSRAMILoll := "0000000000";
CHTOLSRAMOiolL := "0000000000";
CHTOLSRAMlioLL := "0000000000";
CHTOLSRAMiiOLL := "0000000000";
CHTOLSRAMO0oll := "0000000000";
CHTOLSRAML0Oll := "0000000000";
CHTOLSRAMi0oLL := "0000000000";
CHTOLSRAMo1OLl := "0000000000";
CHTOLSRAML1Oll := "0000000000";
CHTOLSRAMI1oll := "0000000000";
CHTOLSRAMOollL := "0000000000";
CHTOLSRAMLollL := "0000000000";
CHTOLSRAMiolLL := "0000000000";
CHTOLSRAMolLLL := "0000000000";
CHTOLSRAMlLLll := "0000000000";
CHTOLSRAMiLLll := "0000000000";
CHTOLSRAMOILll := "0000000000";
CHTOLSRAMlILLl := "0000000000";
CHTOLSRAMIILll := "0000000000";
CHTOLSRAMO0lll := "0000000000";
CHTOLSRAML0lLL := "0000000000";
CHTOLSRAMi0LLL := "0000000000";
CHTOLSRAMO1lll := "0000000000";
CHTOLSRAML1Lll := "0000000000";
CHTOLSRAMI1Lll := "0000000000";
CHTOLSRAMOOill := "0000000000";
CHTOLSRAMloiLL := "0000000000";
CHTOLSRAMiOILl := "0000000000";
CHTOLSRAMOLill := "0000000000";
CHTOLSRAMLLill := "00";
CHTOLSRAMiLILl := "00";
CHTOLSRAMLlilL := "11";
CHTOLSRAMIlilL := "11";
case uSRam_NUM_loCAtioNS_dwIDth32 is
when 128 =>
CHTOLSRAMIIl0 := "011";
CHTOLSRAMi11OL := CHTOLSRAMOl1(6 downto 0)&"000";
CHTOLSRAMiOLll := CHTOLSRAMll1(6 downto 0)&"000";
CHTOLSRAMI00ol := "0000000000"&CHTOLSRAMlO1(7 downto 0);
CHTOLSRAMOIlol := wen;
CHTOLSRAMoiILL := CHTOLSRAMo0LI(7 downto 0);
when 256 =>
CHTOLSRAMO0l0 := "010";
CHTOLSRAMiIL0 := "010";
CHTOLSRAMOOoll := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAMi11OL := CHTOLSRAMol1(7 downto 0)&"00";
CHTOLSRAMOLllL := CHTOLSRAMll1(7 downto 0)&"00";
CHTOLSRAMIollL := CHTOLSRAMll1(7 downto 0)&"00";
CHTOLSRAMO10ol := "00000000000000"&CHTOLSRAMlo1(7 downto 4);
CHTOLSRAMi00OL := "00000000000000"&CHTOLSRAMlo1(3 downto 0);
CHTOLSRAMLiloL := Wen;
CHTOLSRAMOiloL := Wen;
CHTOLSRAMOIill := CHTOLSRAML0lI(3 downto 0)&CHTOLSRAMO0li(3 downto 0);
when 384 =>
CHTOLSRAML0l0 := "010";
CHTOLSRAMO0L0 := "010";
CHTOLSRAMIIl0 := "011";
CHTOLSRAMloOLL := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAMOoolL := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAMI11ol := CHTOLSRAMoL1(6 downto 0)&"000";
CHTOLSRAMLLllL := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMOllLL := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMIOlll := CHTOLSRAMLL1(6 downto 0)&"000";
CHTOLSRAMl10Ol := "00000000000000"&CHTOLSRAMlo1(7 downto 4);
CHTOLSRAMo10OL := "00000000000000"&CHTOLSRAMLO1(3 downto 0);
CHTOLSRAMI00ol := "0000000000"&CHTOLSRAMlo1(7 downto 0);
case CHTOLSRAMoL1(8 downto 6) is
when "000"
| "001"
| "010"
| "011" =>
CHTOLSRAMIIlol := Wen;
CHTOLSRAMliLOl := wen;
CHTOLSRAMoILOl := '0';
when "100"
| "101" =>
CHTOLSRAMIILol := '0';
CHTOLSRAMLiloL := '0';
CHTOLSRAMoILOl := WEn;
when others =>
CHTOLSRAMIiloL := '0';
CHTOLSRAMliLOl := '0';
CHTOLSRAMOIlol := '0';
end case;
case CHTOLSRAMl1Ll(8 downto 6) is
when "000"
| "001"
| "010"
| "011" =>
CHTOLSRAMoiiLL := CHTOLSRAMI0Li(3 downto 0)&CHTOLSRAMl0LI(3 downto 0);
when "100"
| "101" =>
CHTOLSRAMoIILl := CHTOLSRAMo0LI(7 downto 0);
when others =>
CHTOLSRAMOiilL := ( others => '0');
end case;
when 512 =>
CHTOLSRAMI0l0 := "001";
CHTOLSRAMl0L0 := "001";
CHTOLSRAMo0l0 := "001";
CHTOLSRAMIIl0 := "001";
CHTOLSRAMIOOll := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMlOOLl := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMoooLL := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAMI11OL := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAMILlll := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMLLlll := CHTOLSRAMLl1(8 downto 0)&'0';
CHTOLSRAMOllLL := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMIOllL := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMI10ol := "0000000000000000"&CHTOLSRAMlO1(7 downto 6);
CHTOLSRAML10ol := "0000000000000000"&CHTOLSRAMLo1(5 downto 4);
CHTOLSRAMo10Ol := "0000000000000000"&CHTOLSRAMLO1(3 downto 2);
CHTOLSRAMI00ol := "0000000000000000"&CHTOLSRAMLO1(1 downto 0);
CHTOLSRAMo0LOl := wEN;
CHTOLSRAMiILOl := wen;
CHTOLSRAMlilOL := Wen;
CHTOLSRAMOIloL := wEN;
CHTOLSRAMoiiLL := CHTOLSRAMO1li(1 downto 0)&CHTOLSRAMI0li(1 downto 0)&CHTOLSRAMl0LI(1 downto 0)&CHTOLSRAMO0li(1 downto 0);
when 640 =>
CHTOLSRAMi0L0 := "001";
CHTOLSRAML0L0 := "001";
CHTOLSRAMO0l0 := "001";
CHTOLSRAMiIL0 := "001";
CHTOLSRAMliL0 := "011";
CHTOLSRAMioOLL := CHTOLSRAMOl1(8 downto 0)&'0';
CHTOLSRAMLoolL := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAMOoolL := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMI11OL := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMl11OL := CHTOLSRAMOl1(6 downto 0)&"000";
CHTOLSRAMILllL := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMlllLL := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMOLLll := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMioLLL := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMloLLL := CHTOLSRAMlL1(6 downto 0)&"000";
CHTOLSRAMI10oL := "0000000000000000"&CHTOLSRAMLo1(7 downto 6);
CHTOLSRAMl10Ol := "0000000000000000"&CHTOLSRAMLO1(5 downto 4);
CHTOLSRAMO10oL := "0000000000000000"&CHTOLSRAMLO1(3 downto 2);
CHTOLSRAMi00OL := "0000000000000000"&CHTOLSRAMLo1(1 downto 0);
CHTOLSRAML00ol := "0000000000"&CHTOLSRAMLO1(7 downto 0);
case CHTOLSRAMOL1(9 downto 6) is
when "0000"
| "0001"
| "0010"
| "0011"
| "0100"
| "0101"
| "0110"
| "0111" =>
CHTOLSRAMO0lol := WEN;
CHTOLSRAMIiloL := weN;
CHTOLSRAMLIlol := Wen;
CHTOLSRAMoiLOL := wEN;
CHTOLSRAMILlol := '0';
when "1000"
| "1001" =>
CHTOLSRAMo0lOL := '0';
CHTOLSRAMiiLOL := '0';
CHTOLSRAMliLOL := '0';
CHTOLSRAMoiLOL := '0';
CHTOLSRAMiLLOl := WEN;
when others =>
CHTOLSRAMo0LOL := '0';
CHTOLSRAMiiLOL := '0';
CHTOLSRAMLIlol := '0';
CHTOLSRAMoiLOl := '0';
CHTOLSRAMIllOL := '0';
end case;
case CHTOLSRAML1Ll(9 downto 6) is
when "0000"
| "0001"
| "0010"
| "0011"
| "0100"
| "0101"
| "0110"
| "0111" =>
CHTOLSRAMOIilL := CHTOLSRAMo1LI(1 downto 0)&CHTOLSRAMI0li(1 downto 0)&CHTOLSRAML0li(1 downto 0)&CHTOLSRAMO0Li(1 downto 0);
when "1000"
| "1001" =>
CHTOLSRAMOiilL := CHTOLSRAMiiLI(7 downto 0);
when others =>
CHTOLSRAMOIill := ( others => '0');
end case;
when 768 =>
CHTOLSRAMO1L0 := "001";
CHTOLSRAMI0l0 := "001";
CHTOLSRAML0L0 := "001";
CHTOLSRAMo0L0 := "001";
CHTOLSRAMiIL0 := "010";
CHTOLSRAMlIL0 := "010";
CHTOLSRAMolOLl := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMiOOLl := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAMLOoll := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAMoooLL := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMI11oL := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAMl11Ol := CHTOLSRAMOl1(7 downto 0)&"00";
CHTOLSRAMoiLLL := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMillLL := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMLLlll := CHTOLSRAMLl1(8 downto 0)&'0';
CHTOLSRAMOLllL := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMiOLLl := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMlolLL := CHTOLSRAMlL1(7 downto 0)&"00";
CHTOLSRAMoO1Ol := "0000000000000000"&CHTOLSRAMLo1(7 downto 6);
CHTOLSRAMI10ol := "0000000000000000"&CHTOLSRAMlo1(5 downto 4);
CHTOLSRAMl10Ol := "0000000000000000"&CHTOLSRAMLO1(3 downto 2);
CHTOLSRAMO10ol := "0000000000000000"&CHTOLSRAMLo1(1 downto 0);
CHTOLSRAMi00OL := "00000000000000"&CHTOLSRAMLo1(7 downto 4);
CHTOLSRAML00ol := "00000000000000"&CHTOLSRAMlo1(3 downto 0);
case CHTOLSRAMOL1(9 downto 6) is
when "0000"
| "0001"
| "0010"
| "0011"
| "0100"
| "0101"
| "0110"
| "0111" =>
CHTOLSRAMl0LOl := weN;
CHTOLSRAMO0lol := weN;
CHTOLSRAMIIlol := weN;
CHTOLSRAMLILol := WEn;
CHTOLSRAMoiLOL := '0';
CHTOLSRAMILloL := '0';
when "1000"
| "1001"
| "1010"
| "1011" =>
CHTOLSRAML0Lol := '0';
CHTOLSRAMO0lol := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMLiloL := '0';
CHTOLSRAMoILOl := wEN;
CHTOLSRAMILlol := Wen;
when others =>
CHTOLSRAMl0LOL := '0';
CHTOLSRAMo0LOL := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMlilOL := '0';
CHTOLSRAMOILol := '0';
CHTOLSRAMILloL := '0';
end case;
case CHTOLSRAML1ll(9 downto 6) is
when "0000"
| "0001"
| "0010"
| "0011"
| "0100"
| "0101"
| "0110"
| "0111" =>
CHTOLSRAMoiiLL := CHTOLSRAML1li(1 downto 0)&CHTOLSRAMo1lI(1 downto 0)&CHTOLSRAMi0LI(1 downto 0)&CHTOLSRAML0li(1 downto 0);
when "1000"
| "1001"
| "1010"
| "1011" =>
CHTOLSRAMoIILl := CHTOLSRAMO0li(3 downto 0)&CHTOLSRAMIILi(3 downto 0);
when others =>
CHTOLSRAMOIill := ( others => '0');
end case;
when 896 =>
CHTOLSRAML1l0 := "001";
CHTOLSRAMo1l0 := "001";
CHTOLSRAMi0L0 := "001";
CHTOLSRAML0l0 := "001";
CHTOLSRAMo0L0 := "010";
CHTOLSRAMIil0 := "010";
CHTOLSRAMLil0 := "011";
CHTOLSRAMLloLL := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAMolOLl := CHTOLSRAMOl1(8 downto 0)&'0';
CHTOLSRAMIOoll := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMloOLl := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMooOLL := CHTOLSRAMoL1(7 downto 0)&"00";
CHTOLSRAMI11ol := CHTOLSRAMol1(7 downto 0)&"00";
CHTOLSRAMl11OL := CHTOLSRAMol1(6 downto 0)&"000";
CHTOLSRAMliLLl := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMOIllL := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMILLll := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMLlllL := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMOllLL := CHTOLSRAMll1(7 downto 0)&"00";
CHTOLSRAMIOLll := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMlolLL := CHTOLSRAMll1(6 downto 0)&"000";
CHTOLSRAMLo1OL := "0000000000000000"&CHTOLSRAMLo1(7 downto 6);
CHTOLSRAMoO1Ol := "0000000000000000"&CHTOLSRAMLO1(5 downto 4);
CHTOLSRAMI10oL := "0000000000000000"&CHTOLSRAMLO1(3 downto 2);
CHTOLSRAMl10OL := "0000000000000000"&CHTOLSRAMlo1(1 downto 0);
CHTOLSRAMO10oL := "00000000000000"&CHTOLSRAMLO1(7 downto 4);
CHTOLSRAMI00OL := "00000000000000"&CHTOLSRAMlo1(3 downto 0);
CHTOLSRAMl00OL := "0000000000"&CHTOLSRAMlo1(7 downto 0);
case CHTOLSRAMOl1(9 downto 6) is
when "0000"
| "0001"
| "0010"
| "0011"
| "0100"
| "0101"
| "0110"
| "0111" =>
CHTOLSRAMI0lol := WEn;
CHTOLSRAMl0lOL := wen;
CHTOLSRAMo0Lol := wEN;
CHTOLSRAMIiloL := WEn;
CHTOLSRAMlilOL := '0';
CHTOLSRAMoilOL := '0';
CHTOLSRAMillOL := '0';
when "1000"
| "1001"
| "1010"
| "1011" =>
CHTOLSRAMI0lol := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIILol := '0';
CHTOLSRAMLiloL := Wen;
CHTOLSRAMoiLOL := weN;
CHTOLSRAMILlol := '0';
when "1100"
| "1101" =>
CHTOLSRAMI0lOL := '0';
CHTOLSRAML0lOL := '0';
CHTOLSRAMo0lOL := '0';
CHTOLSRAMiilOL := '0';
CHTOLSRAMlilOL := '0';
CHTOLSRAMoilOL := '0';
CHTOLSRAMILlol := WEn;
when others =>
CHTOLSRAMI0lol := '0';
CHTOLSRAML0loL := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMiiLOl := '0';
CHTOLSRAMLIlol := '0';
CHTOLSRAMoiLOl := '0';
CHTOLSRAMILloL := '0';
end case;
case CHTOLSRAMl1LL(9 downto 6) is
when "0000"
| "0001"
| "0010"
| "0011"
| "0100"
| "0101"
| "0110"
| "0111" =>
CHTOLSRAMOiilL := CHTOLSRAMI1li(1 downto 0)&CHTOLSRAMl1LI(1 downto 0)&CHTOLSRAMO1li(1 downto 0)&CHTOLSRAMI0li(1 downto 0);
when "1000"
| "1001"
| "1010"
| "1011" =>
CHTOLSRAMOIIll := CHTOLSRAML0Li(3 downto 0)&CHTOLSRAMO0li(3 downto 0);
when "1100"
| "1101" =>
CHTOLSRAMoiiLL := CHTOLSRAMiILI(7 downto 0);
when others =>
CHTOLSRAMoIIll := ( others => '0');
end case;
when 1024 =>
CHTOLSRAMI1l0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMo1L0 := "000";
CHTOLSRAMi0L0 := "000";
CHTOLSRAMl0l0 := "000";
CHTOLSRAMO0L0 := "000";
CHTOLSRAMiIL0 := "000";
CHTOLSRAMlil0 := "000";
CHTOLSRAMILOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLLoll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMolOLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMIOolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMlOOLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMoOOLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMi11Ol := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMl11OL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMiILLl := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMlilLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMoiLLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMillLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMLlllL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMOLlll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMiolLL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMLOLll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMiO1ol := "00000000000000000"&CHTOLSRAMLo1(7);
CHTOLSRAMLO1ol := "00000000000000000"&CHTOLSRAMLO1(6);
CHTOLSRAMoo1OL := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMI10oL := "00000000000000000"&CHTOLSRAMLo1(4);
CHTOLSRAML10OL := "00000000000000000"&CHTOLSRAMlO1(3);
CHTOLSRAMo10Ol := "00000000000000000"&CHTOLSRAMLO1(2);
CHTOLSRAMI00oL := "00000000000000000"&CHTOLSRAMlo1(1);
CHTOLSRAML00oL := "00000000000000000"&CHTOLSRAMlO1(0);
CHTOLSRAMo1LOl := WEN;
CHTOLSRAMI0lol := Wen;
CHTOLSRAMl0LOL := weN;
CHTOLSRAMo0Lol := weN;
CHTOLSRAMiILOl := Wen;
CHTOLSRAMlilOL := wen;
CHTOLSRAMOiloL := WEN;
CHTOLSRAMILLol := wEN;
CHTOLSRAMoiiLL := CHTOLSRAMoOII(0)&CHTOLSRAMI1li(0)&CHTOLSRAML1lI(0)&CHTOLSRAMO1li(0)&CHTOLSRAMI0li(0)&CHTOLSRAMl0lI(0)&CHTOLSRAMO0lI(0)&CHTOLSRAMIILi(0);
when 1152 =>
CHTOLSRAMOOi0 := "000";
CHTOLSRAMI1l0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMo1l0 := "000";
CHTOLSRAMi0L0 := "000";
CHTOLSRAML0l0 := "000";
CHTOLSRAMO0l0 := "000";
CHTOLSRAMiil0 := "000";
CHTOLSRAMlIL0 := "011";
CHTOLSRAMOIoll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMIlolL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMLlolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMoLOLl := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMIOoll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLoolL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMOoolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMi11OL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAML11oL := CHTOLSRAMoL1(6 downto 0)&"000";
CHTOLSRAMo0LLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMiILll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMlilLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMoILll := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMIllLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMLLLll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMollLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMIOlll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMlolLL := CHTOLSRAMlL1(6 downto 0)&"000";
CHTOLSRAMol1OL := "00000000000000000"&CHTOLSRAMlO1(7);
CHTOLSRAMiO1Ol := "00000000000000000"&CHTOLSRAMlO1(6);
CHTOLSRAMLO1oL := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMOO1oL := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMi10ol := "00000000000000000"&CHTOLSRAMLo1(3);
CHTOLSRAML10oL := "00000000000000000"&CHTOLSRAMlO1(2);
CHTOLSRAMo10Ol := "00000000000000000"&CHTOLSRAMLo1(1);
CHTOLSRAMi00OL := "00000000000000000"&CHTOLSRAMLO1(0);
CHTOLSRAMl00Ol := "0000000000"&CHTOLSRAMlO1(7 downto 0);
case CHTOLSRAMol1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMl1LOl := WEn;
CHTOLSRAMO1loL := wen;
CHTOLSRAMi0LOL := weN;
CHTOLSRAMl0Lol := wEN;
CHTOLSRAMO0Lol := weN;
CHTOLSRAMIILol := WEn;
CHTOLSRAMLiloL := wen;
CHTOLSRAMoiLOL := wen;
CHTOLSRAMilLOL := '0';
when "10000"
| "10001" =>
CHTOLSRAML1Lol := '0';
CHTOLSRAMO1loL := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAML0lOL := '0';
CHTOLSRAMo0LOL := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMLIlol := '0';
CHTOLSRAMoILol := '0';
CHTOLSRAMiLLol := WEn;
when others =>
CHTOLSRAML1loL := '0';
CHTOLSRAMo1LOl := '0';
CHTOLSRAMI0Lol := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMo0lOL := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMLILol := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMilLOL := '0';
end case;
case CHTOLSRAMl1lL(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMoiiLL := CHTOLSRAMloiI(0)&CHTOLSRAMOOii(0)&CHTOLSRAMi1LI(0)&CHTOLSRAML1Li(0)&CHTOLSRAMO1li(0)&CHTOLSRAMI0Li(0)&CHTOLSRAML0Li(0)&CHTOLSRAMO0Li(0);
when "10000"
| "10001" =>
CHTOLSRAMoiILL := CHTOLSRAMiILI(7 downto 0);
when others =>
CHTOLSRAMOIIll := ( others => '0');
end case;
when 1280 =>
CHTOLSRAMloi0 := "000";
CHTOLSRAMOoi0 := "000";
CHTOLSRAMi1L0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMO1L0 := "000";
CHTOLSRAMI0L0 := "000";
CHTOLSRAML0l0 := "000";
CHTOLSRAMo0L0 := "000";
CHTOLSRAMIIL0 := "010";
CHTOLSRAMLIl0 := "010";
CHTOLSRAMLIOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMoIOLl := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMiLOLl := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLLoll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMoloLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMIoolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMlOOll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMOOOll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMi11Ol := CHTOLSRAMol1(7 downto 0)&"00";
CHTOLSRAML11oL := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAML0lll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMO0lll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMIILll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMlILll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMoILLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMILLll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMLlllL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMoLLLl := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMIOlll := CHTOLSRAMLl1(7 downto 0)&"00";
CHTOLSRAMLOlll := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMLL1ol := "00000000000000000"&CHTOLSRAMLo1(7);
CHTOLSRAMOl1OL := "00000000000000000"&CHTOLSRAMLO1(6);
CHTOLSRAMIO1ol := "00000000000000000"&CHTOLSRAMlO1(5);
CHTOLSRAMlO1Ol := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMoO1ol := "00000000000000000"&CHTOLSRAMlo1(3);
CHTOLSRAMI10ol := "00000000000000000"&CHTOLSRAMLo1(2);
CHTOLSRAMl10ol := "00000000000000000"&CHTOLSRAMLo1(1);
CHTOLSRAMO10ol := "00000000000000000"&CHTOLSRAMLO1(0);
CHTOLSRAMI00ol := "00000000000000"&CHTOLSRAMlO1(7 downto 4);
CHTOLSRAMl00Ol := "00000000000000"&CHTOLSRAMLO1(3 downto 0);
case CHTOLSRAMOl1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMi1lOL := Wen;
CHTOLSRAMl1LOL := wEN;
CHTOLSRAMO1lol := wen;
CHTOLSRAMi0LOL := weN;
CHTOLSRAML0Lol := WEn;
CHTOLSRAMO0loL := wen;
CHTOLSRAMiILOl := wEN;
CHTOLSRAMlILOl := Wen;
CHTOLSRAMoiLOL := '0';
CHTOLSRAMILlol := '0';
when "10000"
| "10001"
| "10010"
| "10011" =>
CHTOLSRAMi1LOL := '0';
CHTOLSRAMl1LOl := '0';
CHTOLSRAMO1Lol := '0';
CHTOLSRAMi0Lol := '0';
CHTOLSRAMl0Lol := '0';
CHTOLSRAMO0loL := '0';
CHTOLSRAMiILOl := '0';
CHTOLSRAMLIlol := '0';
CHTOLSRAMoiLOL := WEn;
CHTOLSRAMillOL := wen;
when others =>
CHTOLSRAMi1LOL := '0';
CHTOLSRAML1lol := '0';
CHTOLSRAMo1lOL := '0';
CHTOLSRAMI0Lol := '0';
CHTOLSRAML0loL := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIILol := '0';
CHTOLSRAMLIlol := '0';
CHTOLSRAMoiLOL := '0';
CHTOLSRAMiLLol := '0';
end case;
case CHTOLSRAML1ll(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMoiiLL := CHTOLSRAMIOIi(0)&CHTOLSRAMLOii(0)&CHTOLSRAMooII(0)&CHTOLSRAMi1LI(0)&CHTOLSRAMl1lI(0)&CHTOLSRAMO1li(0)&CHTOLSRAMi0LI(0)&CHTOLSRAMl0LI(0);
when "10000"
| "10001"
| "10010"
| "10011" =>
CHTOLSRAMoiiLL := CHTOLSRAMo0LI(3 downto 0)&CHTOLSRAMiilI(3 downto 0);
when others =>
CHTOLSRAMOIill := ( others => '0');
end case;
when 1408 =>
CHTOLSRAMIoi0 := "000";
CHTOLSRAMLoi0 := "000";
CHTOLSRAMooI0 := "000";
CHTOLSRAMi1l0 := "000";
CHTOLSRAMl1L0 := "000";
CHTOLSRAMO1L0 := "000";
CHTOLSRAMi0L0 := "000";
CHTOLSRAML0L0 := "000";
CHTOLSRAMO0l0 := "010";
CHTOLSRAMiiL0 := "010";
CHTOLSRAMLIl0 := "011";
CHTOLSRAMIIOll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMLiolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMoiOLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMiLOLl := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMLLOll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMoloLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMioOLl := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMLoolL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMOOoll := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAMI11OL := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAML11ol := CHTOLSRAMOL1(6 downto 0)&"000";
CHTOLSRAMi0LLl := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMl0LLl := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMO0lLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMiilLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMLIlll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMoILll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMilLLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMllLLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMoLLLl := CHTOLSRAMll1(7 downto 0)&"00";
CHTOLSRAMiOLLl := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMlOLLl := CHTOLSRAMLL1(6 downto 0)&"000";
CHTOLSRAMil1OL := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMlL1Ol := "00000000000000000"&CHTOLSRAMLO1(6);
CHTOLSRAMoL1Ol := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMiO1ol := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMLO1ol := "00000000000000000"&CHTOLSRAMlo1(3);
CHTOLSRAMoO1Ol := "00000000000000000"&CHTOLSRAMlo1(2);
CHTOLSRAMI10oL := "00000000000000000"&CHTOLSRAMLO1(1);
CHTOLSRAMl10Ol := "00000000000000000"&CHTOLSRAMLO1(0);
CHTOLSRAMO10ol := "00000000000000"&CHTOLSRAMlO1(7 downto 4);
CHTOLSRAMi00Ol := "00000000000000"&CHTOLSRAMLO1(3 downto 0);
CHTOLSRAML00OL := "0000000000"&CHTOLSRAMLO1(7 downto 0);
case CHTOLSRAMol1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMOoiOL := WEn;
CHTOLSRAMI1loL := Wen;
CHTOLSRAML1lol := WEn;
CHTOLSRAMO1loL := wEN;
CHTOLSRAMI0lol := weN;
CHTOLSRAMl0LOL := WEn;
CHTOLSRAMO0loL := Wen;
CHTOLSRAMiilOL := weN;
CHTOLSRAMlILol := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMiLLOl := '0';
when "10000"
| "10001"
| "10010"
| "10011" =>
CHTOLSRAMOOioL := '0';
CHTOLSRAMi1LOL := '0';
CHTOLSRAMl1LOL := '0';
CHTOLSRAMo1LOL := '0';
CHTOLSRAMi0lOL := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMO0lol := '0';
CHTOLSRAMiILOl := '0';
CHTOLSRAMLIlol := wEN;
CHTOLSRAMOILol := WEN;
CHTOLSRAMiLLOl := '0';
when "10100"
| "10101" =>
CHTOLSRAMoOIol := '0';
CHTOLSRAMI1loL := '0';
CHTOLSRAML1loL := '0';
CHTOLSRAMo1LOl := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAML0lol := '0';
CHTOLSRAMO0lol := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMLILol := '0';
CHTOLSRAMoILOl := '0';
CHTOLSRAMILLol := wen;
when others =>
CHTOLSRAMOoioL := '0';
CHTOLSRAMi1Lol := '0';
CHTOLSRAMl1LOl := '0';
CHTOLSRAMo1LOL := '0';
CHTOLSRAMI0loL := '0';
CHTOLSRAMl0lOL := '0';
CHTOLSRAMO0lol := '0';
CHTOLSRAMiILOl := '0';
CHTOLSRAMLILol := '0';
CHTOLSRAMoilOL := '0';
CHTOLSRAMILlol := '0';
end case;
case CHTOLSRAML1ll(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMOIIll := CHTOLSRAMoliI(0)&CHTOLSRAMIoii(0)&CHTOLSRAMlOII(0)&CHTOLSRAMooiI(0)&CHTOLSRAMi1LI(0)&CHTOLSRAMl1lI(0)&CHTOLSRAMo1lI(0)&CHTOLSRAMi0LI(0);
when "10000"
| "10001"
| "10010"
| "10011" =>
CHTOLSRAMOIIll := CHTOLSRAMl0LI(3 downto 0)&CHTOLSRAMo0lI(3 downto 0);
when "10100"
| "10101" =>
CHTOLSRAMOIill := CHTOLSRAMiiLI(7 downto 0);
when others =>
CHTOLSRAMoIILl := ( others => '0');
end case;
when 1536 =>
CHTOLSRAMoli0 := "000";
CHTOLSRAMioI0 := "000";
CHTOLSRAMLoi0 := "000";
CHTOLSRAMoOI0 := "000";
CHTOLSRAMI1L0 := "000";
CHTOLSRAMl1l0 := "000";
CHTOLSRAMO1l0 := "000";
CHTOLSRAMI0l0 := "000";
CHTOLSRAMl0l0 := "001";
CHTOLSRAMo0l0 := "001";
CHTOLSRAMIIl0 := "001";
CHTOLSRAMlil0 := "001";
CHTOLSRAMo0OLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMiioLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMLIolL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMOiolL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMiLOLl := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMlloLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMOlolL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMIOolL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLOOll := CHTOLSRAMOl1(8 downto 0)&'0';
CHTOLSRAMooOLl := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMI11ol := CHTOLSRAMoL1(8 downto 0)&'0';
CHTOLSRAML11oL := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMo1Lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMI0Lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAML0llL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMO0lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMIIlll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMlILll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMoILLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMiLLLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMllLLL := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMOlllL := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMIollL := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMlOLLl := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMOI1oL := "00000000000000000"&CHTOLSRAMlO1(7);
CHTOLSRAMil1Ol := "00000000000000000"&CHTOLSRAMLo1(6);
CHTOLSRAMLl1OL := "00000000000000000"&CHTOLSRAMlo1(5);
CHTOLSRAMOL1ol := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMio1OL := "00000000000000000"&CHTOLSRAMlO1(3);
CHTOLSRAMlO1ol := "00000000000000000"&CHTOLSRAMLo1(2);
CHTOLSRAMoo1OL := "00000000000000000"&CHTOLSRAMlo1(1);
CHTOLSRAMi10Ol := "00000000000000000"&CHTOLSRAMLo1(0);
CHTOLSRAMl10OL := "0000000000000000"&CHTOLSRAMLO1(7 downto 6);
CHTOLSRAMo10Ol := "0000000000000000"&CHTOLSRAMlo1(5 downto 4);
CHTOLSRAMi00OL := "0000000000000000"&CHTOLSRAMLO1(3 downto 2);
CHTOLSRAML00ol := "0000000000000000"&CHTOLSRAMLo1(1 downto 0);
case CHTOLSRAMol1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMloiOL := WEN;
CHTOLSRAMOoiOL := weN;
CHTOLSRAMI1lol := wen;
CHTOLSRAML1Lol := weN;
CHTOLSRAMO1lol := wen;
CHTOLSRAMi0LOL := wEN;
CHTOLSRAML0loL := wen;
CHTOLSRAMo0Lol := wEN;
CHTOLSRAMiILol := '0';
CHTOLSRAMliLOl := '0';
CHTOLSRAMoilOL := '0';
CHTOLSRAMIlloL := '0';
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMLOIol := '0';
CHTOLSRAMoOIOl := '0';
CHTOLSRAMI1lol := '0';
CHTOLSRAMl1LOL := '0';
CHTOLSRAMO1loL := '0';
CHTOLSRAMI0loL := '0';
CHTOLSRAML0loL := '0';
CHTOLSRAMo0lOL := '0';
CHTOLSRAMIIlol := wen;
CHTOLSRAMlilOL := wEN;
CHTOLSRAMOILol := WEn;
CHTOLSRAMIlloL := weN;
when others =>
CHTOLSRAMlOIOl := '0';
CHTOLSRAMOoiOL := '0';
CHTOLSRAMi1Lol := '0';
CHTOLSRAML1loL := '0';
CHTOLSRAMO1lOL := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAML0Lol := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMlILol := '0';
CHTOLSRAMoiLOl := '0';
CHTOLSRAMIlloL := '0';
end case;
case CHTOLSRAMl1LL(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMoIILl := CHTOLSRAMLliI(0)&CHTOLSRAMoLIi(0)&CHTOLSRAMIOii(0)&CHTOLSRAMloII(0)&CHTOLSRAMoOIi(0)&CHTOLSRAMI1Li(0)&CHTOLSRAMl1LI(0)&CHTOLSRAMo1lI(0);
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMOiilL := CHTOLSRAMI0li(1 downto 0)&CHTOLSRAML0Li(1 downto 0)&CHTOLSRAMO0li(1 downto 0)&CHTOLSRAMIIli(1 downto 0);
when others =>
CHTOLSRAMOiiLL := ( others => '0');
end case;
when 1664 =>
CHTOLSRAMllI0 := "000";
CHTOLSRAMOli0 := "000";
CHTOLSRAMIOi0 := "000";
CHTOLSRAMlOI0 := "000";
CHTOLSRAMOOi0 := "000";
CHTOLSRAMI1l0 := "000";
CHTOLSRAMl1L0 := "000";
CHTOLSRAMO1l0 := "000";
CHTOLSRAMi0L0 := "001";
CHTOLSRAMl0l0 := "001";
CHTOLSRAMO0l0 := "001";
CHTOLSRAMIil0 := "001";
CHTOLSRAMlIL0 := "011";
CHTOLSRAML0oll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMo0OLl := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMiIOLl := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMLiolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMOIOll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMiLOLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMLLOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMOLolL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMiOOLl := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMLOolL := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMOOoll := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMI11oL := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMl11OL := CHTOLSRAMOL1(6 downto 0)&"000";
CHTOLSRAML1llL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMo1LLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMI0lLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMl0LLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMO0lll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMIILll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMliLLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMoILLl := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMiLLll := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMlLLLl := CHTOLSRAMlL1(8 downto 0)&'0';
CHTOLSRAMolLLL := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMIOLll := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMLollL := CHTOLSRAMll1(6 downto 0)&"000";
CHTOLSRAMlI1ol := "00000000000000000"&CHTOLSRAMlO1(7);
CHTOLSRAMoI1Ol := "00000000000000000"&CHTOLSRAMLO1(6);
CHTOLSRAMIL1ol := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMll1OL := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMoL1Ol := "00000000000000000"&CHTOLSRAMLO1(3);
CHTOLSRAMIO1ol := "00000000000000000"&CHTOLSRAMlo1(2);
CHTOLSRAMLO1ol := "00000000000000000"&CHTOLSRAMlo1(1);
CHTOLSRAMoo1OL := "00000000000000000"&CHTOLSRAMLo1(0);
CHTOLSRAMi10OL := "0000000000000000"&CHTOLSRAMlo1(7 downto 6);
CHTOLSRAMl10Ol := "0000000000000000"&CHTOLSRAMlo1(5 downto 4);
CHTOLSRAMO10oL := "0000000000000000"&CHTOLSRAMLo1(3 downto 2);
CHTOLSRAMI00ol := "0000000000000000"&CHTOLSRAMlO1(1 downto 0);
CHTOLSRAML00ol := "0000000000"&CHTOLSRAMLo1(7 downto 0);
case CHTOLSRAMOL1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMioiOL := WEn;
CHTOLSRAMlOIOl := WEn;
CHTOLSRAMooIOL := WEn;
CHTOLSRAMI1loL := weN;
CHTOLSRAML1Lol := Wen;
CHTOLSRAMo1LOl := WEn;
CHTOLSRAMi0lOL := Wen;
CHTOLSRAMl0LOL := WEN;
CHTOLSRAMo0Lol := '0';
CHTOLSRAMIilOL := '0';
CHTOLSRAMlILOl := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMIllOL := '0';
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMIoiOL := '0';
CHTOLSRAMloiOL := '0';
CHTOLSRAMoOIol := '0';
CHTOLSRAMI1loL := '0';
CHTOLSRAMl1LOl := '0';
CHTOLSRAMO1lol := '0';
CHTOLSRAMI0Lol := '0';
CHTOLSRAML0lol := '0';
CHTOLSRAMO0lOL := WEn;
CHTOLSRAMIiloL := weN;
CHTOLSRAMliLOL := WEN;
CHTOLSRAMOILol := wEN;
CHTOLSRAMilLOl := '0';
when "11000"
| "11001" =>
CHTOLSRAMioiOL := '0';
CHTOLSRAMLOIol := '0';
CHTOLSRAMOoioL := '0';
CHTOLSRAMI1Lol := '0';
CHTOLSRAML1lOL := '0';
CHTOLSRAMO1lol := '0';
CHTOLSRAMI0lol := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMo0Lol := '0';
CHTOLSRAMiiLOl := '0';
CHTOLSRAMliLOL := '0';
CHTOLSRAMoILol := '0';
CHTOLSRAMilLOl := WEn;
when others =>
CHTOLSRAMIoioL := '0';
CHTOLSRAMLOiol := '0';
CHTOLSRAMOOIol := '0';
CHTOLSRAMi1LOL := '0';
CHTOLSRAML1Lol := '0';
CHTOLSRAMO1loL := '0';
CHTOLSRAMI0lol := '0';
CHTOLSRAML0loL := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIIloL := '0';
CHTOLSRAMlILOl := '0';
CHTOLSRAMoilOL := '0';
CHTOLSRAMILlol := '0';
end case;
case CHTOLSRAML1ll(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMoIIll := CHTOLSRAMILIi(0)&CHTOLSRAMllII(0)&CHTOLSRAMolII(0)&CHTOLSRAMIOii(0)&CHTOLSRAMLOii(0)&CHTOLSRAMooII(0)&CHTOLSRAMi1LI(0)&CHTOLSRAMl1LI(0);
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMOIill := CHTOLSRAMo1lI(1 downto 0)&CHTOLSRAMi0LI(1 downto 0)&CHTOLSRAML0li(1 downto 0)&CHTOLSRAMo0LI(1 downto 0);
when "11000"
| "11001" =>
CHTOLSRAMoIILl := CHTOLSRAMiiLI(7 downto 0);
when others =>
CHTOLSRAMOIill := ( others => '0');
end case;
when 1792 =>
CHTOLSRAMili0 := "000";
CHTOLSRAMlLI0 := "000";
CHTOLSRAMoLI0 := "000";
CHTOLSRAMioi0 := "000";
CHTOLSRAMLOI0 := "000";
CHTOLSRAMOoi0 := "000";
CHTOLSRAMi1l0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMo1L0 := "001";
CHTOLSRAMi0L0 := "001";
CHTOLSRAMl0L0 := "001";
CHTOLSRAMO0L0 := "001";
CHTOLSRAMIil0 := "010";
CHTOLSRAMLIL0 := "010";
CHTOLSRAMI0oll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMl0oLL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMo0OLL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMIIOll := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMliOLl := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMOIolL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMILOll := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMlLOll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMolOLL := CHTOLSRAMOl1(8 downto 0)&'0';
CHTOLSRAMIOoll := CHTOLSRAMOl1(8 downto 0)&'0';
CHTOLSRAMlOOLl := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMOOoll := CHTOLSRAMOl1(8 downto 0)&'0';
CHTOLSRAMi11Ol := CHTOLSRAMoL1(7 downto 0)&"00";
CHTOLSRAMl11OL := CHTOLSRAMOl1(7 downto 0)&"00";
CHTOLSRAMi1lLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMl1LlL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMo1lLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMI0lll := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAML0Lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMo0LLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMIillL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMlILLl := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMoILLl := CHTOLSRAMLl1(8 downto 0)&'0';
CHTOLSRAMILLll := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMLLLll := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMollLL := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMIOlll := CHTOLSRAMLL1(7 downto 0)&"00";
CHTOLSRAMLOlll := CHTOLSRAMLl1(7 downto 0)&"00";
CHTOLSRAMii1Ol := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMLI1ol := "00000000000000000"&CHTOLSRAMlo1(6);
CHTOLSRAMOi1OL := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMil1Ol := "00000000000000000"&CHTOLSRAMLO1(4);
CHTOLSRAMLl1oL := "00000000000000000"&CHTOLSRAMlO1(3);
CHTOLSRAMOL1ol := "00000000000000000"&CHTOLSRAMlo1(2);
CHTOLSRAMiO1Ol := "00000000000000000"&CHTOLSRAMlO1(1);
CHTOLSRAMLO1ol := "00000000000000000"&CHTOLSRAMLo1(0);
CHTOLSRAMOo1oL := "0000000000000000"&CHTOLSRAMLo1(7 downto 6);
CHTOLSRAMI10ol := "0000000000000000"&CHTOLSRAMLO1(5 downto 4);
CHTOLSRAML10oL := "0000000000000000"&CHTOLSRAMLo1(3 downto 2);
CHTOLSRAMO10ol := "0000000000000000"&CHTOLSRAMlo1(1 downto 0);
CHTOLSRAMi00Ol := "00000000000000"&CHTOLSRAMLO1(7 downto 4);
CHTOLSRAML00ol := "00000000000000"&CHTOLSRAMLO1(3 downto 0);
case CHTOLSRAMOL1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMOLiol := weN;
CHTOLSRAMIOioL := weN;
CHTOLSRAMLoiOL := weN;
CHTOLSRAMooIOl := weN;
CHTOLSRAMI1Lol := wen;
CHTOLSRAMl1Lol := Wen;
CHTOLSRAMO1lOL := weN;
CHTOLSRAMI0lol := WEn;
CHTOLSRAML0lOL := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIIlol := '0';
CHTOLSRAMLiloL := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMIlloL := '0';
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMOLIol := '0';
CHTOLSRAMioIOL := '0';
CHTOLSRAMloiOL := '0';
CHTOLSRAMooiOL := '0';
CHTOLSRAMI1loL := '0';
CHTOLSRAML1lol := '0';
CHTOLSRAMO1lOL := '0';
CHTOLSRAMI0lol := '0';
CHTOLSRAML0lOL := wEN;
CHTOLSRAMO0Lol := wEN;
CHTOLSRAMIIlol := WEN;
CHTOLSRAMLIlol := WEN;
CHTOLSRAMOIlol := '0';
CHTOLSRAMILlol := '0';
when "11000"
| "11001"
| "11010"
| "11011" =>
CHTOLSRAMOlioL := '0';
CHTOLSRAMiOIol := '0';
CHTOLSRAMLOiol := '0';
CHTOLSRAMOoioL := '0';
CHTOLSRAMI1lOL := '0';
CHTOLSRAML1lOL := '0';
CHTOLSRAMO1lol := '0';
CHTOLSRAMI0lOL := '0';
CHTOLSRAML0lol := '0';
CHTOLSRAMo0LOL := '0';
CHTOLSRAMiiLOL := '0';
CHTOLSRAMliLOL := '0';
CHTOLSRAMoiLOL := WEn;
CHTOLSRAMIlloL := weN;
when others =>
CHTOLSRAMoliOL := '0';
CHTOLSRAMioIOL := '0';
CHTOLSRAMloIOL := '0';
CHTOLSRAMOOioL := '0';
CHTOLSRAMi1LOl := '0';
CHTOLSRAMl1lOL := '0';
CHTOLSRAMO1loL := '0';
CHTOLSRAMI0loL := '0';
CHTOLSRAML0lol := '0';
CHTOLSRAMO0Lol := '0';
CHTOLSRAMiILol := '0';
CHTOLSRAMlilOL := '0';
CHTOLSRAMoiLOL := '0';
CHTOLSRAMillOL := '0';
end case;
case CHTOLSRAML1lL(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMoiILL := CHTOLSRAMoIII(0)&CHTOLSRAMILIi(0)&CHTOLSRAMLliI(0)&CHTOLSRAMoliI(0)&CHTOLSRAMIOii(0)&CHTOLSRAMlOII(0)&CHTOLSRAMooII(0)&CHTOLSRAMI1li(0);
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMOiilL := CHTOLSRAML1li(1 downto 0)&CHTOLSRAMO1li(1 downto 0)&CHTOLSRAMI0li(1 downto 0)&CHTOLSRAML0li(1 downto 0);
when "11000"
| "11001"
| "11010"
| "11011" =>
CHTOLSRAMoiILL := CHTOLSRAMO0li(3 downto 0)&CHTOLSRAMiILi(3 downto 0);
when others =>
CHTOLSRAMOIilL := ( others => '0');
end case;
when 1920 =>
CHTOLSRAMoII0 := "000";
CHTOLSRAMiLI0 := "000";
CHTOLSRAMllI0 := "000";
CHTOLSRAMOLi0 := "000";
CHTOLSRAMioI0 := "000";
CHTOLSRAMLOI0 := "000";
CHTOLSRAMOOI0 := "000";
CHTOLSRAMi1l0 := "000";
CHTOLSRAML1l0 := "001";
CHTOLSRAMO1L0 := "001";
CHTOLSRAMI0l0 := "001";
CHTOLSRAMl0l0 := "001";
CHTOLSRAMO0l0 := "010";
CHTOLSRAMIIL0 := "010";
CHTOLSRAMliL0 := "011";
CHTOLSRAMO1oll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMI0olL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAML0oLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMO0oll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMIIoll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMLIOll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMOIOll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMiloLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMlLOLl := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMoLOLl := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMioOLL := CHTOLSRAMOL1(8 downto 0)&'0';
CHTOLSRAMlOOLl := CHTOLSRAMol1(8 downto 0)&'0';
CHTOLSRAMOOOll := CHTOLSRAMoL1(7 downto 0)&"00";
CHTOLSRAMi11OL := CHTOLSRAMoL1(7 downto 0)&"00";
CHTOLSRAML11ol := CHTOLSRAMOL1(6 downto 0)&"000";
CHTOLSRAMooiLL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMI1lLL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAML1lll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMO1lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMI0lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMl0LLl := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMo0LLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMIillL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMlILll := CHTOLSRAMLl1(8 downto 0)&'0';
CHTOLSRAMOIllL := CHTOLSRAMll1(8 downto 0)&'0';
CHTOLSRAMILLll := CHTOLSRAMLl1(8 downto 0)&'0';
CHTOLSRAMLLLll := CHTOLSRAMLL1(8 downto 0)&'0';
CHTOLSRAMolLLL := CHTOLSRAMlL1(7 downto 0)&"00";
CHTOLSRAMIOllL := CHTOLSRAMll1(7 downto 0)&"00";
CHTOLSRAMLOLll := CHTOLSRAMLL1(6 downto 0)&"000";
CHTOLSRAMo01ol := "00000000000000000"&CHTOLSRAMlO1(7);
CHTOLSRAMii1OL := "00000000000000000"&CHTOLSRAMLo1(6);
CHTOLSRAMlI1Ol := "00000000000000000"&CHTOLSRAMlO1(5);
CHTOLSRAMOi1OL := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMIL1ol := "00000000000000000"&CHTOLSRAMLO1(3);
CHTOLSRAMll1OL := "00000000000000000"&CHTOLSRAMLO1(2);
CHTOLSRAMol1OL := "00000000000000000"&CHTOLSRAMLo1(1);
CHTOLSRAMiO1Ol := "00000000000000000"&CHTOLSRAMlO1(0);
CHTOLSRAMLO1ol := "0000000000000000"&CHTOLSRAMlO1(7 downto 6);
CHTOLSRAMoo1OL := "0000000000000000"&CHTOLSRAMlO1(5 downto 4);
CHTOLSRAMi10OL := "0000000000000000"&CHTOLSRAMlO1(3 downto 2);
CHTOLSRAMl10Ol := "0000000000000000"&CHTOLSRAMLo1(1 downto 0);
CHTOLSRAMo10OL := "00000000000000"&CHTOLSRAMLO1(7 downto 4);
CHTOLSRAMI00OL := "00000000000000"&CHTOLSRAMLO1(3 downto 0);
CHTOLSRAMl00ol := "0000000000"&CHTOLSRAMLO1(7 downto 0);
case CHTOLSRAMOL1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMLLIol := wEN;
CHTOLSRAMOLiol := Wen;
CHTOLSRAMiOIOl := WEn;
CHTOLSRAMloiOL := Wen;
CHTOLSRAMoOIOl := wEN;
CHTOLSRAMI1loL := Wen;
CHTOLSRAMl1LOL := wEN;
CHTOLSRAMo1LOl := wEN;
CHTOLSRAMI0loL := '0';
CHTOLSRAML0Lol := '0';
CHTOLSRAMO0loL := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMlILOl := '0';
CHTOLSRAMOIlol := '0';
CHTOLSRAMIlloL := '0';
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMlliOL := '0';
CHTOLSRAMolIOL := '0';
CHTOLSRAMiOIOl := '0';
CHTOLSRAMLOIol := '0';
CHTOLSRAMOOiol := '0';
CHTOLSRAMI1Lol := '0';
CHTOLSRAML1lOL := '0';
CHTOLSRAMo1LOl := '0';
CHTOLSRAMi0LOl := weN;
CHTOLSRAMl0LOl := weN;
CHTOLSRAMo0LOl := weN;
CHTOLSRAMIILol := Wen;
CHTOLSRAMliLOl := '0';
CHTOLSRAMoILol := '0';
CHTOLSRAMILLol := '0';
when "11000"
| "11001"
| "11010"
| "11011" =>
CHTOLSRAMLLIol := '0';
CHTOLSRAMolIOl := '0';
CHTOLSRAMIOIol := '0';
CHTOLSRAMlOIOl := '0';
CHTOLSRAMOOIol := '0';
CHTOLSRAMI1Lol := '0';
CHTOLSRAML1loL := '0';
CHTOLSRAMO1loL := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAMl0lOL := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIIlol := '0';
CHTOLSRAMlILOl := Wen;
CHTOLSRAMoiLOL := weN;
CHTOLSRAMILlol := '0';
when "11100"
| "11101" =>
CHTOLSRAMllIOL := '0';
CHTOLSRAMoLIol := '0';
CHTOLSRAMiOIOl := '0';
CHTOLSRAMLOIol := '0';
CHTOLSRAMOOioL := '0';
CHTOLSRAMI1Lol := '0';
CHTOLSRAML1lol := '0';
CHTOLSRAMo1lOL := '0';
CHTOLSRAMi0lOL := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMO0loL := '0';
CHTOLSRAMiilOL := '0';
CHTOLSRAMLIlol := '0';
CHTOLSRAMoiLOl := '0';
CHTOLSRAMILloL := wen;
when others =>
CHTOLSRAMLlioL := '0';
CHTOLSRAMoLIOl := '0';
CHTOLSRAMiOIOl := '0';
CHTOLSRAMLoioL := '0';
CHTOLSRAMooIOL := '0';
CHTOLSRAMi1lOL := '0';
CHTOLSRAML1loL := '0';
CHTOLSRAMo1Lol := '0';
CHTOLSRAMi0LOL := '0';
CHTOLSRAML0lol := '0';
CHTOLSRAMo0Lol := '0';
CHTOLSRAMIIlol := '0';
CHTOLSRAMLIloL := '0';
CHTOLSRAMOILol := '0';
CHTOLSRAMillOL := '0';
end case;
case CHTOLSRAML1ll(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMoiILL := CHTOLSRAMlIII(0)&CHTOLSRAMoIII(0)&CHTOLSRAMIlii(0)&CHTOLSRAMLliI(0)&CHTOLSRAMoLII(0)&CHTOLSRAMIOIi(0)&CHTOLSRAMloII(0)&CHTOLSRAMOOIi(0);
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111" =>
CHTOLSRAMoiiLL := CHTOLSRAMi1LI(1 downto 0)&CHTOLSRAML1li(1 downto 0)&CHTOLSRAMO1li(1 downto 0)&CHTOLSRAMi0Li(1 downto 0);
when "11000"
| "11001"
| "11010"
| "11011" =>
CHTOLSRAMOIIll := CHTOLSRAML0li(3 downto 0)&CHTOLSRAMO0li(3 downto 0);
when "11100"
| "11101" =>
CHTOLSRAMoiILL := CHTOLSRAMIIli(7 downto 0);
when others =>
CHTOLSRAMoIIll := ( others => '0');
end case;
when 2048 =>
CHTOLSRAMLII0 := "000";
CHTOLSRAMOIi0 := "000";
CHTOLSRAMILI0 := "000";
CHTOLSRAMlLI0 := "000";
CHTOLSRAMoli0 := "000";
CHTOLSRAMIOI0 := "000";
CHTOLSRAMlOI0 := "000";
CHTOLSRAMOOI0 := "000";
CHTOLSRAMi1L0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMO1L0 := "000";
CHTOLSRAMi0L0 := "000";
CHTOLSRAML0l0 := "000";
CHTOLSRAMo0L0 := "000";
CHTOLSRAMIIL0 := "000";
CHTOLSRAMliL0 := "000";
CHTOLSRAML1Oll := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMO1oll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMI0olL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAML0olL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMO0oLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMIiolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMlIOLl := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMOIolL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMIloLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLLOll := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMoLOLl := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMIOOll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMLOoll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMoooLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMi11Ol := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMl11ol := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMLOill := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMOOill := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMi1LLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMl1LLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMo1LLl := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMi0LLl := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMl0LLl := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMO0llL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMiiLLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMLILll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMOillL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMillLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMlLLLl := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMolLLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMIOllL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMLOLll := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMl01Ol := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMO01oL := "00000000000000000"&CHTOLSRAMLO1(6);
CHTOLSRAMIi1oL := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMLI1ol := "00000000000000000"&CHTOLSRAMLO1(4);
CHTOLSRAMoi1OL := "00000000000000000"&CHTOLSRAMlo1(3);
CHTOLSRAMiL1Ol := "00000000000000000"&CHTOLSRAMLo1(2);
CHTOLSRAMll1OL := "00000000000000000"&CHTOLSRAMLO1(1);
CHTOLSRAMol1Ol := "00000000000000000"&CHTOLSRAMLo1(0);
CHTOLSRAMio1OL := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMlO1Ol := "00000000000000000"&CHTOLSRAMlo1(6);
CHTOLSRAMoo1OL := "00000000000000000"&CHTOLSRAMLO1(5);
CHTOLSRAMi10Ol := "00000000000000000"&CHTOLSRAMlO1(4);
CHTOLSRAML10oL := "00000000000000000"&CHTOLSRAMLO1(3);
CHTOLSRAMO10oL := "00000000000000000"&CHTOLSRAMlo1(2);
CHTOLSRAMI00oL := "00000000000000000"&CHTOLSRAMlo1(1);
CHTOLSRAMl00ol := "00000000000000000"&CHTOLSRAMLO1(0);
case CHTOLSRAMOl1(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMIliOL := WEN;
CHTOLSRAMlLIOl := WEn;
CHTOLSRAMOlioL := Wen;
CHTOLSRAMioIOl := Wen;
CHTOLSRAMLOIol := Wen;
CHTOLSRAMOOiol := Wen;
CHTOLSRAMI1Lol := weN;
CHTOLSRAML1loL := wEN;
CHTOLSRAMO1lol := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAMl0LOl := '0';
CHTOLSRAMO0lOL := '0';
CHTOLSRAMiILOl := '0';
CHTOLSRAMlILOl := '0';
CHTOLSRAMOilOL := '0';
CHTOLSRAMILloL := '0';
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111"
| "11000"
| "11001"
| "11010"
| "11011"
| "11100"
| "11101"
| "11110"
| "11111" =>
CHTOLSRAMIliOL := '0';
CHTOLSRAMLLioL := '0';
CHTOLSRAMoliOL := '0';
CHTOLSRAMioiOL := '0';
CHTOLSRAMloIOl := '0';
CHTOLSRAMOOIol := '0';
CHTOLSRAMI1loL := '0';
CHTOLSRAML1Lol := '0';
CHTOLSRAMO1loL := weN;
CHTOLSRAMI0Lol := wEN;
CHTOLSRAML0Lol := WEn;
CHTOLSRAMO0loL := Wen;
CHTOLSRAMIiloL := Wen;
CHTOLSRAMLiloL := wen;
CHTOLSRAMOILol := WEn;
CHTOLSRAMillOL := wen;
when others =>
CHTOLSRAMILiol := '0';
CHTOLSRAMLlioL := '0';
CHTOLSRAMOLioL := '0';
CHTOLSRAMIOiol := '0';
CHTOLSRAMLOiol := '0';
CHTOLSRAMOoioL := '0';
CHTOLSRAMI1Lol := '0';
CHTOLSRAML1lol := '0';
CHTOLSRAMO1Lol := '0';
CHTOLSRAMI0lol := '0';
CHTOLSRAML0lol := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIIlol := '0';
CHTOLSRAMLILol := '0';
CHTOLSRAMOILol := '0';
CHTOLSRAMIlloL := '0';
end case;
case CHTOLSRAMl1lL(10 downto 6) is
when "00000"
| "00001"
| "00010"
| "00011"
| "00100"
| "00101"
| "00110"
| "00111"
| "01000"
| "01001"
| "01010"
| "01011"
| "01100"
| "01101"
| "01110"
| "01111" =>
CHTOLSRAMOiilL := CHTOLSRAMiiiI(0)&CHTOLSRAMliII(0)&CHTOLSRAMOIii(0)&CHTOLSRAMiLII(0)&CHTOLSRAMLliI(0)&CHTOLSRAMoLIi(0)&CHTOLSRAMIOii(0)&CHTOLSRAMLoii(0);
when "10000"
| "10001"
| "10010"
| "10011"
| "10100"
| "10101"
| "10110"
| "10111"
| "11000"
| "11001"
| "11010"
| "11011"
| "11100"
| "11101"
| "11110"
| "11111" =>
CHTOLSRAMoIIll := CHTOLSRAMooII(0)&CHTOLSRAMi1LI(0)&CHTOLSRAML1li(0)&CHTOLSRAMo1LI(0)&CHTOLSRAMi0LI(0)&CHTOLSRAML0li(0)&CHTOLSRAMo0LI(0)&CHTOLSRAMiilI(0);
when others =>
CHTOLSRAMOIilL := ( others => '0');
end case;
when 2176 =>
CHTOLSRAMIIi0 := "000";
CHTOLSRAMLIi0 := "000";
CHTOLSRAMOii0 := "000";
CHTOLSRAMIli0 := "000";
CHTOLSRAMlli0 := "000";
CHTOLSRAMoLI0 := "000";
CHTOLSRAMiOI0 := "000";
CHTOLSRAMLOi0 := "000";
CHTOLSRAMoOI0 := "000";
CHTOLSRAMi1L0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMo1L0 := "000";
CHTOLSRAMI0l0 := "000";
CHTOLSRAMl0L0 := "000";
CHTOLSRAMo0l0 := "000";
CHTOLSRAMIil0 := "000";
CHTOLSRAMlil0 := "011";
CHTOLSRAMI1Oll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMl1oLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMo1oLL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMi0OLL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMl0oLL := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMO0oLL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMIIOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLIOll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMOIoll := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMiLOLl := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMLLoll := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMoLOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMiOOLl := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMLOoll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMoOOLl := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMi11OL := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMl11Ol := CHTOLSRAMol1(6 downto 0)&"000";
CHTOLSRAMIoiLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMLOilL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMooiLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMI1llL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMl1Lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMO1lll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMi0LLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAML0llL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMO0lll := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMiiLLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMlilLL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMoiLLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMilLLL := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMLLllL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMOlllL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMiOLLl := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMLOLll := CHTOLSRAMLL1(6 downto 0)&"000";
CHTOLSRAMI01OL := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMl01OL := "00000000000000000"&CHTOLSRAMLO1(6);
CHTOLSRAMO01ol := "00000000000000000"&CHTOLSRAMlO1(5);
CHTOLSRAMIi1oL := "00000000000000000"&CHTOLSRAMlo1(4);
CHTOLSRAMlI1ol := "00000000000000000"&CHTOLSRAMLO1(3);
CHTOLSRAMOi1OL := "00000000000000000"&CHTOLSRAMlo1(2);
CHTOLSRAMIl1oL := "00000000000000000"&CHTOLSRAMLo1(1);
CHTOLSRAMlL1Ol := "00000000000000000"&CHTOLSRAMlo1(0);
CHTOLSRAMOl1oL := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMIo1oL := "00000000000000000"&CHTOLSRAMlO1(6);
CHTOLSRAMlo1OL := "00000000000000000"&CHTOLSRAMlO1(5);
CHTOLSRAMoo1OL := "00000000000000000"&CHTOLSRAMlO1(4);
CHTOLSRAMI10OL := "00000000000000000"&CHTOLSRAMlo1(3);
CHTOLSRAML10ol := "00000000000000000"&CHTOLSRAMlO1(2);
CHTOLSRAMO10oL := "00000000000000000"&CHTOLSRAMLO1(1);
CHTOLSRAMi00OL := "00000000000000000"&CHTOLSRAMlO1(0);
CHTOLSRAML00oL := "0000000000"&CHTOLSRAMlO1(7 downto 0);
case CHTOLSRAMOL1(11 downto 6) is
when "000000"
| "000001"
| "000010"
| "000011"
| "000100"
| "000101"
| "000110"
| "000111"
| "001000"
| "001001"
| "001010"
| "001011"
| "001100"
| "001101"
| "001110"
| "001111" =>
CHTOLSRAMOiioL := wen;
CHTOLSRAMiliOL := weN;
CHTOLSRAMLLiol := wen;
CHTOLSRAMoLIol := WEn;
CHTOLSRAMioiOL := weN;
CHTOLSRAMloiOL := Wen;
CHTOLSRAMOOIol := WEn;
CHTOLSRAMI1Lol := Wen;
CHTOLSRAMl1lOL := '0';
CHTOLSRAMo1lOL := '0';
CHTOLSRAMI0Lol := '0';
CHTOLSRAML0lOL := '0';
CHTOLSRAMo0LOl := '0';
CHTOLSRAMIiloL := '0';
CHTOLSRAMlILol := '0';
CHTOLSRAMOIloL := '0';
CHTOLSRAMILlol := '0';
when "010000"
| "010001"
| "010010"
| "010011"
| "010100"
| "010101"
| "010110"
| "010111"
| "011000"
| "011001"
| "011010"
| "011011"
| "011100"
| "011101"
| "011110"
| "011111" =>
CHTOLSRAMoiiOL := '0';
CHTOLSRAMiliOL := '0';
CHTOLSRAMlLIOl := '0';
CHTOLSRAMOLioL := '0';
CHTOLSRAMiOIOl := '0';
CHTOLSRAMloIOL := '0';
CHTOLSRAMOOIol := '0';
CHTOLSRAMi1LOL := '0';
CHTOLSRAMl1Lol := WEn;
CHTOLSRAMo1LOl := WEn;
CHTOLSRAMi0lOL := Wen;
CHTOLSRAMl0LOl := WEn;
CHTOLSRAMo0lOL := WEN;
CHTOLSRAMIiloL := wEN;
CHTOLSRAMLIloL := WEN;
CHTOLSRAMoilOL := WEn;
CHTOLSRAMIlloL := '0';
when "100000"
| "100001" =>
CHTOLSRAMOiioL := '0';
CHTOLSRAMIliOL := '0';
CHTOLSRAMlliOL := '0';
CHTOLSRAMolIOL := '0';
CHTOLSRAMIOIol := '0';
CHTOLSRAMloIOL := '0';
CHTOLSRAMOOiol := '0';
CHTOLSRAMi1LOl := '0';
CHTOLSRAMl1lOL := '0';
CHTOLSRAMO1loL := '0';
CHTOLSRAMi0LOL := '0';
CHTOLSRAML0loL := '0';
CHTOLSRAMO0lOL := '0';
CHTOLSRAMIilOL := '0';
CHTOLSRAMLiloL := '0';
CHTOLSRAMoilOL := '0';
CHTOLSRAMillOL := WEN;
when others =>
CHTOLSRAMOIioL := '0';
CHTOLSRAMIlioL := '0';
CHTOLSRAMlLIol := '0';
CHTOLSRAMoLIol := '0';
CHTOLSRAMIoioL := '0';
CHTOLSRAMLOIol := '0';
CHTOLSRAMooIOl := '0';
CHTOLSRAMi1LOl := '0';
CHTOLSRAML1Lol := '0';
CHTOLSRAMo1lOL := '0';
CHTOLSRAMI0lol := '0';
CHTOLSRAMl0LOL := '0';
CHTOLSRAMO0lOL := '0';
CHTOLSRAMiILOl := '0';
CHTOLSRAMliLOL := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMILlol := '0';
end case;
case CHTOLSRAML1Ll(11 downto 6) is
when "000000"
| "000001"
| "000010"
| "000011"
| "000100"
| "000101"
| "000110"
| "000111"
| "001000"
| "001001"
| "001010"
| "001011"
| "001100"
| "001101"
| "001110"
| "001111" =>
CHTOLSRAMOIill := CHTOLSRAMo0iI(0)&CHTOLSRAMiIII(0)&CHTOLSRAMliII(0)&CHTOLSRAMOiii(0)&CHTOLSRAMILIi(0)&CHTOLSRAMlliI(0)&CHTOLSRAMoLIi(0)&CHTOLSRAMIoiI(0);
when "010000"
| "010001"
| "010010"
| "010011"
| "010100"
| "010101"
| "010110"
| "010111"
| "011000"
| "011001"
| "011010"
| "011011"
| "011100"
| "011101"
| "011110"
| "011111" =>
CHTOLSRAMOIill := CHTOLSRAMlOII(0)&CHTOLSRAMOOii(0)&CHTOLSRAMi1LI(0)&CHTOLSRAMl1LI(0)&CHTOLSRAMo1LI(0)&CHTOLSRAMi0LI(0)&CHTOLSRAMl0LI(0)&CHTOLSRAMo0LI(0);
when "100000"
| "100001" =>
CHTOLSRAMoiILL := CHTOLSRAMiiLI(7 downto 0);
when others =>
CHTOLSRAMOIIll := ( others => '0');
end case;
when 2304 =>
CHTOLSRAMO0i0 := "000";
CHTOLSRAMIIi0 := "000";
CHTOLSRAMLii0 := "000";
CHTOLSRAMoII0 := "000";
CHTOLSRAMilI0 := "000";
CHTOLSRAMLLI0 := "000";
CHTOLSRAMOLi0 := "000";
CHTOLSRAMioi0 := "000";
CHTOLSRAMloI0 := "000";
CHTOLSRAMOOi0 := "000";
CHTOLSRAMI1l0 := "000";
CHTOLSRAML1l0 := "000";
CHTOLSRAMO1l0 := "000";
CHTOLSRAMI0l0 := "000";
CHTOLSRAMl0l0 := "000";
CHTOLSRAMo0l0 := "000";
CHTOLSRAMIil0 := "010";
CHTOLSRAMLil0 := "010";
CHTOLSRAMooLLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMI1olL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMl1OLl := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMo1OLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMi0oLL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMl0oLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMo0OLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMiiOLl := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMLIoll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMOiolL := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMiLOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMlloLL := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMOLoll := CHTOLSRAMoL1(9 downto 0);
CHTOLSRAMIOOll := CHTOLSRAMOl1(9 downto 0);
CHTOLSRAMlOOLl := CHTOLSRAMOL1(9 downto 0);
CHTOLSRAMOOOll := CHTOLSRAMol1(9 downto 0);
CHTOLSRAMi11OL := CHTOLSRAMOL1(7 downto 0)&"00";
CHTOLSRAML11ol := CHTOLSRAMoL1(7 downto 0)&"00";
CHTOLSRAMOLIll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMIOill := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMloILl := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMoOIll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMi1LLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMl1LLl := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMo1LLl := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMI0llL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMl0LLL := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMO0llL := CHTOLSRAMLl1(9 downto 0);
CHTOLSRAMIillL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMlILll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMoILLl := CHTOLSRAMLL1(9 downto 0);
CHTOLSRAMIlllL := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMLLlll := CHTOLSRAMlL1(9 downto 0);
CHTOLSRAMOLlll := CHTOLSRAMll1(9 downto 0);
CHTOLSRAMIOLll := CHTOLSRAMLl1(7 downto 0)&"00";
CHTOLSRAMLOlll := CHTOLSRAMlL1(7 downto 0)&"00";
CHTOLSRAMO11OL := "00000000000000000"&CHTOLSRAMLO1(7);
CHTOLSRAMI01ol := "00000000000000000"&CHTOLSRAMlO1(6);
CHTOLSRAMl01OL := "00000000000000000"&CHTOLSRAMLo1(5);
CHTOLSRAMO01ol := "00000000000000000"&CHTOLSRAMLo1(4);
CHTOLSRAMii1OL := "00000000000000000"&CHTOLSRAMlO1(3);
CHTOLSRAMLI1ol := "00000000000000000"&CHTOLSRAMlO1(2);
CHTOLSRAMOI1ol := "00000000000000000"&CHTOLSRAMLO1(1);
CHTOLSRAMIL1ol := "00000000000000000"&CHTOLSRAMlo1(0);
CHTOLSRAMll1OL := "00000000000000000"&CHTOLSRAMLo1(7);
CHTOLSRAMOL1oL := "00000000000000000"&CHTOLSRAMlO1(6);
CHTOLSRAMio1OL := "00000000000000000"&CHTOLSRAMlO1(5);
CHTOLSRAMlo1OL := "00000000000000000"&CHTOLSRAMLO1(4);
CHTOLSRAMoo1OL := "00000000000000000"&CHTOLSRAMLo1(3);
CHTOLSRAMI10oL := "00000000000000000"&CHTOLSRAMlo1(2);
CHTOLSRAML10ol := "00000000000000000"&CHTOLSRAMLO1(1);
CHTOLSRAMO10ol := "00000000000000000"&CHTOLSRAMLO1(0);
CHTOLSRAMi00oL := "00000000000000"&CHTOLSRAMLO1(7 downto 4);
CHTOLSRAML00oL := "00000000000000"&CHTOLSRAMlO1(3 downto 0);
case CHTOLSRAMOL1(11 downto 6) is
when "000000"
| "000001"
| "000010"
| "000011"
| "000100"
| "000101"
| "000110"
| "000111"
| "001000"
| "001001"
| "001010"
| "001011"
| "001100"
| "001101"
| "001110"
| "001111" =>
CHTOLSRAMliIOL := wen;
CHTOLSRAMoiIOL := WEn;
CHTOLSRAMILIol := weN;
CHTOLSRAMlliOL := Wen;
CHTOLSRAMoLIol := WEn;
CHTOLSRAMioIOL := wen;
CHTOLSRAMLOIol := Wen;
CHTOLSRAMOOiol := Wen;
CHTOLSRAMI1Lol := '0';
CHTOLSRAML1lOL := '0';
CHTOLSRAMO1lol := '0';
CHTOLSRAMi0LOl := '0';
CHTOLSRAMl0lOL := '0';
CHTOLSRAMO0loL := '0';
CHTOLSRAMIILol := '0';
CHTOLSRAMLILol := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMillOL := '0';
when "010000"
| "010001"
| "010010"
| "010011"
| "010100"
| "010101"
| "010110"
| "010111"
| "011000"
| "011001"
| "011010"
| "011011"
| "011100"
| "011101"
| "011110"
| "011111" =>
CHTOLSRAMLIiol := '0';
CHTOLSRAMoiiOL := '0';
CHTOLSRAMiliOL := '0';
CHTOLSRAMLLIol := '0';
CHTOLSRAMOlioL := '0';
CHTOLSRAMioIOL := '0';
CHTOLSRAMLOIol := '0';
CHTOLSRAMoOIOl := '0';
CHTOLSRAMI1lol := Wen;
CHTOLSRAML1loL := weN;
CHTOLSRAMo1LOl := WEn;
CHTOLSRAMi0LOL := wEN;
CHTOLSRAML0loL := wen;
CHTOLSRAMO0loL := wen;
CHTOLSRAMIIlol := WEn;
CHTOLSRAMlilOL := WEn;
CHTOLSRAMOilOL := '0';
CHTOLSRAMILLol := '0';
when "100000"
| "100001"
| "100010"
| "100011" =>
CHTOLSRAMlIIOl := '0';
CHTOLSRAMOIioL := '0';
CHTOLSRAMilIOL := '0';
CHTOLSRAMLLiol := '0';
CHTOLSRAMOlioL := '0';
CHTOLSRAMiOIol := '0';
CHTOLSRAMLOIol := '0';
CHTOLSRAMOOiol := '0';
CHTOLSRAMi1lOL := '0';
CHTOLSRAMl1Lol := '0';
CHTOLSRAMo1LOl := '0';
CHTOLSRAMi0Lol := '0';
CHTOLSRAML0loL := '0';
CHTOLSRAMo0lOL := '0';
CHTOLSRAMIILol := '0';
CHTOLSRAMLILol := '0';
CHTOLSRAMOIlol := wEN;
CHTOLSRAMILlol := weN;
when others =>
CHTOLSRAMLIiol := '0';
CHTOLSRAMoIIol := '0';
CHTOLSRAMILioL := '0';
CHTOLSRAMLLioL := '0';
CHTOLSRAMOlioL := '0';
CHTOLSRAMIoiOL := '0';
CHTOLSRAMlOIOl := '0';
CHTOLSRAMooIOL := '0';
CHTOLSRAMI1loL := '0';
CHTOLSRAML1loL := '0';
CHTOLSRAMO1lol := '0';
CHTOLSRAMI0lol := '0';
CHTOLSRAML0Lol := '0';
CHTOLSRAMO0lol := '0';
CHTOLSRAMiILOl := '0';
CHTOLSRAMlILOl := '0';
CHTOLSRAMOiloL := '0';
CHTOLSRAMiLLOl := '0';
end case;
case CHTOLSRAML1ll(11 downto 6) is
when "000000"
| "000001"
| "000010"
| "000011"
| "000100"
| "000101"
| "000110"
| "000111"
| "001000"
| "001001"
| "001010"
| "001011"
| "001100"
| "001101"
| "001110"
| "001111" =>
CHTOLSRAMOIill := CHTOLSRAML0iI(0)&CHTOLSRAMO0ii(0)&CHTOLSRAMIiii(0)&CHTOLSRAMlIIi(0)&CHTOLSRAMoiII(0)&CHTOLSRAMIliI(0)&CHTOLSRAMLLIi(0)&CHTOLSRAMoliI(0);
when "010000"
| "010001"
| "010010"
| "010011"
| "010100"
| "010101"
| "010110"
| "010111"
| "011000"
| "011001"
| "011010"
| "011011"
| "011100"
| "011101"
| "011110"
| "011111" =>
CHTOLSRAMoIILl := CHTOLSRAMIoii(0)&CHTOLSRAMLoii(0)&CHTOLSRAMOOIi(0)&CHTOLSRAMI1li(0)&CHTOLSRAMl1LI(0)&CHTOLSRAMo1LI(0)&CHTOLSRAMi0LI(0)&CHTOLSRAMl0LI(0);
when "100000"
| "100001"
| "100010"
| "100011" =>
CHTOLSRAMoiILL := CHTOLSRAMo0LI(3 downto 0)&CHTOLSRAMIILi(3 downto 0);
when others =>
CHTOLSRAMoIILl := ( others => '0');
end case;
when others =>
null
;
end case;
wIDTh0 <= CHTOLSRAMLil0;
WidtH1 <= CHTOLSRAMIIl0;
wiDTh2 <= CHTOLSRAMo0L0;
CHTOLSRAMI1ll <= CHTOLSRAMl0L0;
CHTOLSRAMooIL <= CHTOLSRAMi0L0;
CHTOLSRAMLoil <= CHTOLSRAMO1l0;
CHTOLSRAMIoil <= CHTOLSRAMl1l0;
CHTOLSRAMolIL <= CHTOLSRAMi1L0;
CHTOLSRAMllIL <= CHTOLSRAMooI0;
CHTOLSRAMILil <= CHTOLSRAMlOI0;
CHTOLSRAMoiIL <= CHTOLSRAMioi0;
CHTOLSRAMLiil <= CHTOLSRAMOLi0;
CHTOLSRAMiIIL <= CHTOLSRAMllI0;
CHTOLSRAMo0iL <= CHTOLSRAMILi0;
CHTOLSRAML0Il <= CHTOLSRAMoii0;
CHTOLSRAMI0il <= CHTOLSRAMlII0;
CHTOLSRAMo1iL <= CHTOLSRAMIIi0;
CHTOLSRAMl1IL <= CHTOLSRAMO0i0;
CHTOLSRAMi1IL <= CHTOLSRAMillOL;
CHTOLSRAMOO0l <= CHTOLSRAMoiLOL;
CHTOLSRAMlo0L <= CHTOLSRAMlilOL;
CHTOLSRAMIo0l <= CHTOLSRAMIILol;
CHTOLSRAMoL0l <= CHTOLSRAMo0lOL;
CHTOLSRAMLl0l <= CHTOLSRAML0lol;
CHTOLSRAMiL0l <= CHTOLSRAMi0lOL;
CHTOLSRAMOi0l <= CHTOLSRAMo1LOl;
CHTOLSRAMli0L <= CHTOLSRAML1loL;
CHTOLSRAMIi0l <= CHTOLSRAMi1LOl;
CHTOLSRAMo00L <= CHTOLSRAMOoioL;
CHTOLSRAMl00L <= CHTOLSRAMlOIOl;
CHTOLSRAMi00L <= CHTOLSRAMIoioL;
CHTOLSRAMO10l <= CHTOLSRAMoliOL;
CHTOLSRAML10l <= CHTOLSRAMLLIol;
CHTOLSRAMI10l <= CHTOLSRAMiLIOl;
CHTOLSRAMoo1L <= CHTOLSRAMOIiol;
CHTOLSRAMLO1l <= CHTOLSRAMliIOl;
CHTOLSRAMIo1l <= CHTOLSRAMIIioL;
CHTOLSRAMOl1l <= CHTOLSRAMO0Iol;
CHTOLSRAMLL1l <= CHTOLSRAMl0IOL;
CHTOLSRAMil1L <= CHTOLSRAMI0ioL;
CHTOLSRAMOi1l <= CHTOLSRAMO1Iol;
CHTOLSRAMlI1L <= CHTOLSRAML1ioL;
CHTOLSRAMII1l <= CHTOLSRAMi1iOL;
CHTOLSRAMo01L <= CHTOLSRAMoo0Ol;
CHTOLSRAMl01L <= CHTOLSRAMlo0OL;
CHTOLSRAMI01l <= CHTOLSRAMiO0ol;
CHTOLSRAMo11L <= CHTOLSRAMol0Ol;
CHTOLSRAMl11L <= CHTOLSRAMll0OL;
CHTOLSRAMI11l <= CHTOLSRAMIL0ol;
CHTOLSRAMOOoi <= CHTOLSRAMOI0ol;
CHTOLSRAMLOoi <= CHTOLSRAMlI0ol;
CHTOLSRAMioOI <= CHTOLSRAMIi0oL;
CHTOLSRAMOLOi <= CHTOLSRAMo00ol;
CHTOLSRAMILoi <= CHTOLSRAML00oL;
CHTOLSRAMoiOI <= CHTOLSRAMi00Ol;
CHTOLSRAMlIOI <= CHTOLSRAMO10ol;
CHTOLSRAMiIOI <= CHTOLSRAML10oL;
CHTOLSRAMO0oI <= CHTOLSRAMi10OL;
CHTOLSRAMl0OI <= CHTOLSRAMoO1ol;
CHTOLSRAMI0Oi <= CHTOLSRAMLo1oL;
CHTOLSRAMO1oi <= CHTOLSRAMIo1oL;
CHTOLSRAML1oi <= CHTOLSRAMol1OL;
CHTOLSRAMI1Oi <= CHTOLSRAMlL1Ol;
CHTOLSRAMooLI <= CHTOLSRAMiL1ol;
CHTOLSRAMLOli <= CHTOLSRAMoi1Ol;
CHTOLSRAMiOLI <= CHTOLSRAMLi1oL;
CHTOLSRAMOllI <= CHTOLSRAMIi1oL;
CHTOLSRAMLlli <= CHTOLSRAMO01OL;
CHTOLSRAMilLI <= CHTOLSRAML01ol;
CHTOLSRAMoILI <= CHTOLSRAMI01ol;
CHTOLSRAMLili <= CHTOLSRAMo11OL;
CHTOLSRAMi0II <= CHTOLSRAMl11Ol;
CHTOLSRAMo1II <= CHTOLSRAMi11Ol;
CHTOLSRAMl1II <= CHTOLSRAMoOOll;
CHTOLSRAMI1ii <= CHTOLSRAMLoolL;
CHTOLSRAMOO0i <= CHTOLSRAMioOLl;
CHTOLSRAMlo0I <= CHTOLSRAMOLolL;
CHTOLSRAMIo0i <= CHTOLSRAMllOLL;
CHTOLSRAMoL0i <= CHTOLSRAMILoll;
CHTOLSRAMLL0i <= CHTOLSRAMOIOll;
CHTOLSRAMil0I <= CHTOLSRAMlIOLl;
CHTOLSRAMoI0I <= CHTOLSRAMIIOll;
CHTOLSRAMLI0i <= CHTOLSRAMo0Oll;
CHTOLSRAMiI0I <= CHTOLSRAML0olL;
CHTOLSRAMO00i <= CHTOLSRAMI0oLL;
CHTOLSRAMl00I <= CHTOLSRAMO1olL;
CHTOLSRAMI00i <= CHTOLSRAML1oll;
CHTOLSRAMO10i <= CHTOLSRAMi1OLl;
CHTOLSRAML10i <= CHTOLSRAMOOlll;
CHTOLSRAMI10i <= CHTOLSRAMloLLL;
CHTOLSRAMoo1I <= CHTOLSRAMioLLL;
CHTOLSRAMLo1i <= CHTOLSRAMOlllL;
CHTOLSRAMio1I <= CHTOLSRAMlllLL;
CHTOLSRAMOl1I <= CHTOLSRAMillLL;
CHTOLSRAMll1I <= CHTOLSRAMoILLl;
CHTOLSRAMIl1i <= CHTOLSRAMLIlll;
CHTOLSRAMOi1i <= CHTOLSRAMiiLLL;
CHTOLSRAMli1I <= CHTOLSRAMo0LLL;
CHTOLSRAMii1I <= CHTOLSRAMl0lLL;
CHTOLSRAMO01I <= CHTOLSRAMi0Lll;
CHTOLSRAMl01i <= CHTOLSRAMO1llL;
CHTOLSRAMI01i <= CHTOLSRAMl1LLl;
CHTOLSRAMo11I <= CHTOLSRAMi1LLl;
CHTOLSRAMl11I <= CHTOLSRAMooILL;
CHTOLSRAMi11I <= CHTOLSRAMlOILl;
CHTOLSRAMooO0 <= CHTOLSRAMiOILl;
CHTOLSRAMlOO0 <= CHTOLSRAMOLill;
CHTOLSRAMi111 <= CHTOLSRAMLLill;
CHTOLSRAMoooOL <= CHTOLSRAMiliLL;
CHTOLSRAMill0 <= CHTOLSRAMOIIll;
end process;
CHTOLSRAMo0ILl: rAM64x18
port map (A_doUT => CHTOLSRAML0ii,
B_doUT => open ,
a_ADdr_CLk => clk,
B_aDDR_clK => CLK,
a_aDDR_eN => '1',
b_ADdr_EN => '1',
a_aDDr_lAT => '1',
b_ADdr_LAt => '1',
A_addR_arsT_N => CHTOLSRAMiL1,
B_Addr_Arst_N => CHTOLSRAMil1,
a_ADdr_SRSt_n => '1',
b_ADdr_SRst_N => '1',
a_DOut_CLK => '1',
b_dOUT_clK => '1',
A_douT_en => '1',
b_DOut_EN => '1',
A_doUT_lat => '1',
B_DouT_Lat => '1',
A_douT_ArsT_N => CHTOLSRAMIl1,
B_douT_arsT_N => CHTOLSRAMIL1,
A_doUT_srST_n => '1',
B_douT_Srst_N => '1',
a_ADdr => CHTOLSRAMloo0,
b_ADDr => CHTOLSRAMLoo0,
A_WidTH => CHTOLSRAML1il,
B_widTH => CHTOLSRAML1il,
a_Blk => CHTOLSRAMI111,
b_Blk => CHTOLSRAMOoooL,
A_en => '1',
b_eN => '1',
C_clk => clK,
C_AddR => CHTOLSRAML10i,
c_DIn => CHTOLSRAMlilI,
C_weN => CHTOLSRAMlo1L,
C_blK => "11",
C_widTH => CHTOLSRAML1il,
C_En => '1',
Sii_LOCk => '0',
buSY => CHTOLSRAMiOOOl);
CHTOLSRAML0ill: raM64x18
port map (a_DOut => CHTOLSRAMO0Ii,
B_dOUT => open ,
A_addR_Clk => CLk,
B_aDDR_clK => CLK,
A_adDR_en => '1',
b_Addr_EN => '1',
a_aDDr_lAT => '1',
B_aDDR_laT => '1',
a_aDDR_aRST_n => CHTOLSRAMiL1,
b_ADDr_ARSt_n => CHTOLSRAMIL1,
a_Addr_SRst_N => '1',
b_aDDr_sRST_n => '1',
A_doUT_clk => '1',
B_douT_Clk => '1',
a_Dout_EN => '1',
B_doUT_en => '1',
A_doUT_lat => '1',
b_Dout_LAt => '1',
A_douT_ArsT_N => CHTOLSRAMIL1,
b_DOUt_aRST_n => CHTOLSRAMiL1,
a_DOut_SRst_N => '1',
B_doUT_srsT_N => '1',
a_ADdr => CHTOLSRAMOOo0,
b_ADDr => CHTOLSRAMooo0,
A_wiDTH => CHTOLSRAMo1IL,
B_widTH => CHTOLSRAMo1iL,
A_blk => CHTOLSRAMI111,
b_bLK => CHTOLSRAMOoooL,
a_En => '1',
B_eN => '1',
C_clk => cLK,
C_AddR => CHTOLSRAMO10i,
c_DIn => CHTOLSRAMoILI,
C_weN => CHTOLSRAMOO1l,
C_blK => "11",
C_WidtH => CHTOLSRAMo1IL,
C_en => '1',
sii_LOck => '0',
bUSy => CHTOLSRAMlooOL);
CHTOLSRAMI0Ill: RAm64X18
port map (A_douT => CHTOLSRAMiiII,
B_douT => open ,
A_adDR_clk => clK,
B_adDR_clK => clk,
a_aDDr_eN => '1',
B_adDR_en => '1',
a_Addr_LAt => '1',
B_addR_lat => '1',
A_adDR_arST_n => CHTOLSRAMil1,
B_aDDR_arST_n => CHTOLSRAMil1,
A_addR_srsT_N => '1',
b_Addr_SRst_N => '1',
a_DOUt_cLK => '1',
b_dOUt_cLK => '1',
A_douT_En => '1',
b_DOUt_eN => '1',
a_DOUt_LAT => '1',
B_douT_lat => '1',
a_DOut_ARSt_N => CHTOLSRAMIL1,
b_DOUt_ARSt_n => CHTOLSRAMIL1,
a_DOut_SRst_N => '1',
b_DOUt_SRSt_n => '1',
a_Addr => CHTOLSRAMI11i,
b_ADDr => CHTOLSRAMi11I,
A_widTH => CHTOLSRAMi0IL,
B_widTH => CHTOLSRAMI0il,
a_bLK => CHTOLSRAMi111,
b_bLK => CHTOLSRAMOOOol,
a_EN => '1',
B_en => '1',
C_clK => clK,
c_ADDr => CHTOLSRAMi00I,
c_dIN => CHTOLSRAMILli,
c_WEN => CHTOLSRAMI10l,
c_bLK => "11",
c_WIdth => CHTOLSRAMi0IL,
C_en => '1',
sii_Lock => '0',
Busy => CHTOLSRAMolOOL);
CHTOLSRAMO1ilL: RAm64X18
port map (a_DOUt => CHTOLSRAMLiiI,
b_dOUt => open ,
A_Addr_Clk => clK,
B_addR_Clk => cLK,
A_adDR_en => '1',
b_aDDr_eN => '1',
A_addR_Lat => '1',
B_AddR_Lat => '1',
a_ADDr_aRST_n => CHTOLSRAMil1,
B_adDR_arST_n => CHTOLSRAMil1,
A_adDR_srsT_n => '1',
b_ADDr_SRSt_n => '1',
A_douT_Clk => '1',
b_dOUt_cLK => '1',
A_Dout_EN => '1',
b_DOUt_eN => '1',
a_DOUt_lAT => '1',
b_dOUT_laT => '1',
A_douT_ArsT_N => CHTOLSRAMil1,
B_doUT_arsT_n => CHTOLSRAMIl1,
A_doUT_srST_n => '1',
B_Dout_Srst_N => '1',
A_aDDR => CHTOLSRAML11i,
b_Addr => CHTOLSRAMl11I,
A_wiDTh => CHTOLSRAMl0Il,
b_WIDth => CHTOLSRAMl0IL,
A_blK => CHTOLSRAMi111,
B_blK => CHTOLSRAMooOOL,
a_eN => '1',
b_EN => '1',
C_clK => CLK,
c_aDDR => CHTOLSRAMl00i,
c_dIN => CHTOLSRAMllLI,
C_wen => CHTOLSRAML10l,
c_bLK => "11",
C_wiDTH => CHTOLSRAMl0iL,
C_en => '1',
sII_loCK => '0',
busY => CHTOLSRAMLLool);
CHTOLSRAML1Ill: RAm64X18
port map (a_DOUt => CHTOLSRAMOIIi,
B_doUT => open ,
a_aDDR_cLK => clK,
B_Addr_Clk => CLK,
a_aDDR_en => '1',
b_aDDR_eN => '1',
A_addR_Lat => '1',
B_addR_lat => '1',
A_AddR_Arst_N => CHTOLSRAMIl1,
B_addR_arsT_N => CHTOLSRAMIl1,
A_addR_srsT_N => '1',
B_addR_Srst_N => '1',
A_doUT_clk => '1',
b_DOut_CLk => '1',
A_dOUT_en => '1',
B_douT_En => '1',
a_DOut_LAt => '1',
b_DOUt_LAT => '1',
A_dOUT_arST_n => CHTOLSRAMIl1,
b_Dout_ARst_N => CHTOLSRAMIL1,
a_Dout_SRst_N => '1',
B_doUT_srsT_N => '1',
A_adDR => CHTOLSRAMo11I,
b_ADDr => CHTOLSRAMo11i,
a_wIDth => CHTOLSRAMO0Il,
b_WIDth => CHTOLSRAMo0iL,
A_Blk => CHTOLSRAMI111,
b_BLk => CHTOLSRAMOOool,
a_EN => '1',
B_en => '1',
c_CLK => clk,
c_ADdr => CHTOLSRAMO00i,
c_DIN => CHTOLSRAMoLLI,
C_weN => CHTOLSRAMo10L,
C_blK => "11",
C_wiDTH => CHTOLSRAMo0IL,
C_en => '1',
sII_loCK => '0',
Busy => CHTOLSRAMILool);
CHTOLSRAMI1ill: RAm64X18
port map (A_doUT => CHTOLSRAMILii,
B_dOUT => open ,
a_ADdr_CLk => cLK,
B_adDR_clK => Clk,
a_ADDr_eN => '1',
b_ADDr_EN => '1',
A_adDR_laT => '1',
B_addR_Lat => '1',
A_aDDR_arST_n => CHTOLSRAMIL1,
b_Addr_ARst_N => CHTOLSRAMiL1,
a_ADDr_sRSt_n => '1',
b_aDDR_sRST_n => '1',
A_doUT_clk => '1',
B_doUT_clk => '1',
A_douT_en => '1',
b_Dout_EN => '1',
a_DOUt_lAT => '1',
b_DOUt_lAT => '1',
A_doUT_arST_n => CHTOLSRAMil1,
B_douT_Arst_N => CHTOLSRAMIL1,
A_Dout_Srst_N => '1',
b_DOUt_sRSt_n => '1',
a_ADdr => CHTOLSRAMI01i,
b_ADDr => CHTOLSRAMi01I,
a_wIDth => CHTOLSRAMIIil,
b_WIdth => CHTOLSRAMiIIl,
a_bLK => CHTOLSRAMI111,
b_BLk => CHTOLSRAMOooOL,
A_en => '1',
b_EN => '1',
c_CLK => clk,
c_ADDr => CHTOLSRAMii0I,
c_DIN => CHTOLSRAMiOLI,
c_WEN => CHTOLSRAMi00L,
C_blK => "11",
C_widTH => CHTOLSRAMiiiL,
c_eN => '1',
SII_loCK => '0',
Busy => CHTOLSRAMOIooL);
CHTOLSRAMOo0LL: Ram64X18
port map (a_dOUt => CHTOLSRAMLLii,
b_dOUt => open ,
A_addR_clk => CLk,
B_adDR_clK => Clk,
a_ADDr_EN => '1',
B_Addr_En => '1',
a_ADdr_LAt => '1',
B_AddR_Lat => '1',
A_addR_Arst_N => CHTOLSRAMiL1,
b_aDDr_aRST_n => CHTOLSRAMIL1,
a_ADdr_SRst_N => '1',
B_Addr_SRst_N => '1',
A_doUT_clk => '1',
b_dOUt_cLK => '1',
A_doUT_en => '1',
B_DouT_En => '1',
a_DOut_LAT => '1',
b_DOUt_lAT => '1',
A_doUT_arST_n => CHTOLSRAMiL1,
b_dOUt_aRST_n => CHTOLSRAMIL1,
a_DOUt_SRSt_n => '1',
B_doUT_srsT_N => '1',
a_aDDr => CHTOLSRAMl01I,
b_ADdr => CHTOLSRAML01i,
A_WidtH => CHTOLSRAMlIIL,
b_WIDth => CHTOLSRAMLIil,
A_blK => CHTOLSRAMI111,
b_BLk => CHTOLSRAMoOOOl,
a_EN => '1',
B_en => '1',
C_clk => cLK,
c_ADdr => CHTOLSRAMLI0i,
c_dIN => CHTOLSRAMLoli,
C_Wen => CHTOLSRAML00l,
c_BLk => "11",
C_WidTH => CHTOLSRAMLiil,
C_en => '1',
SIi_lOCK => '0',
bUSY => CHTOLSRAMliOOL);
CHTOLSRAMLo0lL: rAM64x18
port map (a_DOut => CHTOLSRAMOlii,
b_DOut => open ,
a_ADdr_CLk => Clk,
b_ADdr_CLk => clK,
A_aDDR_en => '1',
b_ADdr_EN => '1',
a_ADdr_LAT => '1',
b_ADdr_LAt => '1',
a_ADDr_aRSt_n => CHTOLSRAMiL1,
b_ADdr_ARst_N => CHTOLSRAMIL1,
A_AddR_Srst_n => '1',
b_Addr_Srst_N => '1',
a_DOut_CLK => '1',
b_DOUt_cLK => '1',
a_dOUT_eN => '1',
B_douT_En => '1',
A_douT_lat => '1',
b_DOut_LAT => '1',
A_douT_arsT_N => CHTOLSRAMil1,
b_dOUT_arST_n => CHTOLSRAMiL1,
a_DOut_SRSt_n => '1',
b_DOUt_SRSt_n => '1',
A_adDR => CHTOLSRAMo01i,
b_ADdr => CHTOLSRAMO01i,
A_wIDTh => CHTOLSRAMOIIl,
b_wIDth => CHTOLSRAMoiiL,
A_blk => CHTOLSRAMi111,
B_Blk => CHTOLSRAMoOOOl,
a_eN => '1',
b_EN => '1',
c_CLk => clK,
C_Addr => CHTOLSRAMoI0I,
C_diN => CHTOLSRAMoolI,
c_Wen => CHTOLSRAMo00L,
C_blK => "11",
c_WidtH => CHTOLSRAMOiil,
c_EN => '1',
sII_loCK => '0',
Busy => CHTOLSRAMiIOOl);
CHTOLSRAMIO0ll: rAM64x18
port map (a_DOut => CHTOLSRAMIoii,
B_doUT => open ,
a_ADdr_CLk => clk,
b_ADDr_CLK => clk,
a_ADDr_eN => '1',
B_addR_En => '1',
a_ADDr_LAT => '1',
B_adDR_laT => '1',
A_AddR_Arst_N => CHTOLSRAMIl1,
b_ADdr_ARst_N => CHTOLSRAMIl1,
A_AddR_Srst_N => '1',
b_aDDr_sRST_n => '1',
a_DOut_CLk => '1',
B_dOUT_clK => '1',
A_douT_en => '1',
b_DOUt_eN => '1',
A_doUT_lat => '1',
b_DOut_LAt => '1',
a_Dout_ARst_N => CHTOLSRAMIL1,
b_DOUt_ARSt_n => CHTOLSRAMIL1,
a_DOut_SRst_N => '1',
B_doUT_srST_n => '1',
A_adDR => CHTOLSRAMiI1I,
B_adDR => CHTOLSRAMII1i,
a_wIDTh => CHTOLSRAMILIl,
B_wIDTh => CHTOLSRAMILIl,
A_blK => CHTOLSRAMI111,
b_Blk => CHTOLSRAMOoooL,
A_En => '1',
B_En => '1',
C_clK => CLk,
c_ADdr => CHTOLSRAMil0I,
C_diN => CHTOLSRAMi1oI,
C_Wen => CHTOLSRAMII0l,
C_bLK => "11",
C_widTH => CHTOLSRAMiliL,
c_En => '1',
SIi_lOCk => '0',
BusY => CHTOLSRAMO0ool);
CHTOLSRAMOl0LL: Ram64X18
port map (a_DOut => CHTOLSRAMLoii,
B_doUT => open ,
a_ADDr_cLK => clK,
b_ADdr_CLk => cLK,
A_addR_En => '1',
b_ADdr_EN => '1',
a_ADDr_LAT => '1',
b_aDDr_lAT => '1',
a_aDDR_arST_n => CHTOLSRAMiL1,
B_aDDR_arST_n => CHTOLSRAMIL1,
a_aDDr_sRST_n => '1',
B_aDDR_srST_n => '1',
a_DOut_CLK => '1',
B_doUT_clk => '1',
A_dOUT_en => '1',
B_doUT_en => '1',
a_DOUt_LAT => '1',
B_dOUT_laT => '1',
A_douT_ArsT_N => CHTOLSRAMIl1,
b_DOut_ARst_N => CHTOLSRAMIl1,
a_Dout_SRst_N => '1',
B_doUT_srST_n => '1',
A_adDR => CHTOLSRAMLi1I,
b_ADdr => CHTOLSRAMLi1i,
a_WIdtH => CHTOLSRAMllIL,
B_wiDTH => CHTOLSRAMLLIl,
a_bLK => CHTOLSRAMI111,
B_blK => CHTOLSRAMooOOl,
a_EN => '1',
B_en => '1',
c_cLK => Clk,
C_addR => CHTOLSRAMll0I,
C_din => CHTOLSRAML1oI,
C_wen => CHTOLSRAMli0L,
C_blk => "11",
C_wiDTH => CHTOLSRAMlliL,
C_En => '1',
Sii_LOck => '0',
BUSy => CHTOLSRAML0ooL);
CHTOLSRAMLl0LL: Ram64X18
port map (a_DOUt => CHTOLSRAMOOii,
b_DOut => open ,
A_addR_clk => clK,
b_ADdr_CLk => clK,
a_ADdr_EN => '1',
B_aDDR_en => '1',
A_AddR_Lat => '1',
b_ADDr_lAT => '1',
A_adDR_arST_n => CHTOLSRAMiL1,
B_adDR_arST_n => CHTOLSRAMil1,
A_AddR_Srst_N => '1',
B_adDR_srST_n => '1',
a_DOUt_CLK => '1',
b_DOUt_CLK => '1',
a_dOUt_eN => '1',
b_DOut_EN => '1',
a_dOUT_lAT => '1',
B_DouT_Lat => '1',
A_doUT_arST_n => CHTOLSRAMIL1,
b_DOUt_aRSt_n => CHTOLSRAMIL1,
A_Dout_Srst_N => '1',
b_Dout_SRst_N => '1',
a_ADdr => CHTOLSRAMoI1I,
B_adDR => CHTOLSRAMOI1i,
A_wIDTh => CHTOLSRAMolIL,
B_WidTH => CHTOLSRAMOLIl,
a_bLK => CHTOLSRAMi111,
B_blk => CHTOLSRAMoOOOl,
a_eN => '1',
B_En => '1',
C_Clk => clk,
C_aDDR => CHTOLSRAMoL0I,
C_diN => CHTOLSRAMO1Oi,
C_weN => CHTOLSRAMoI0l,
C_blk => "11",
C_wiDTh => CHTOLSRAMOlil,
c_EN => '1',
SII_lOCK => '0',
buSY => CHTOLSRAMI0Ool);
CHTOLSRAMiL0Ll: raM64x18
port map (a_dOUt => CHTOLSRAMI1li,
b_DOUt => open ,
a_ADdr_CLK => clK,
b_ADdr_CLK => Clk,
A_aDDR_en => '1',
b_aDDr_eN => '1',
a_ADdr_LAt => '1',
B_adDR_laT => '1',
a_ADDr_ARSt_n => CHTOLSRAMIL1,
b_Addr_Arst_N => CHTOLSRAMIL1,
a_ADdr_SRSt_N => '1',
B_adDR_srST_n => '1',
a_DOut_CLk => '1',
B_doUT_clk => '1',
a_DOUt_EN => '1',
B_douT_En => '1',
A_dOUT_laT => '1',
b_DOut_LAT => '1',
A_doUT_arsT_n => CHTOLSRAMIL1,
b_DOUt_ARSt_n => CHTOLSRAMiL1,
A_doUT_srST_n => '1',
b_DOut_SRst_N => '1',
a_ADdr => CHTOLSRAMIl1i,
b_ADdr => CHTOLSRAMil1I,
A_WidTH => CHTOLSRAMIOIl,
B_wIDTh => CHTOLSRAMIoil,
a_BLk => CHTOLSRAMI111,
b_BLk => CHTOLSRAMOoooL,
a_En => '1',
B_En => '1',
C_Clk => Clk,
C_adDR => CHTOLSRAMio0I,
c_DIN => CHTOLSRAMI0oI,
c_wEN => CHTOLSRAMIl0L,
c_Blk => "11",
c_WIDth => CHTOLSRAMioIL,
c_En => '1',
SII_loCK => '0',
buSY => CHTOLSRAMo1oOL);
CHTOLSRAMoi0LL: ram64X18
port map (a_DOut => CHTOLSRAMl1lI,
b_dOUt => open ,
a_ADDr_CLK => clk,
b_ADDr_CLK => Clk,
a_aDDr_eN => '1',
B_AddR_En => '1',
A_aDDR_laT => '1',
B_AddR_Lat => '1',
A_AddR_Arst_N => CHTOLSRAMil1,
B_Addr_Arst_N => CHTOLSRAMIl1,
a_ADdr_SRSt_N => '1',
b_Addr_Srst_N => '1',
A_doUT_clK => '1',
b_Dout_CLk => '1',
A_douT_En => '1',
B_doUT_en => '1',
A_Dout_Lat => '1',
B_douT_lat => '1',
a_DOUt_ARSt_n => CHTOLSRAMil1,
B_doUT_arST_n => CHTOLSRAMil1,
A_doUT_srST_n => '1',
b_DOUt_sRSt_n => '1',
a_aDDR => CHTOLSRAMlL1I,
B_adDR => CHTOLSRAMLL1i,
a_wIDTh => CHTOLSRAMlOIL,
B_wIDTh => CHTOLSRAMLOil,
a_bLK => CHTOLSRAMI111,
B_blK => CHTOLSRAMoOOOl,
a_EN => '1',
b_eN => '1',
c_cLK => CLk,
C_addR => CHTOLSRAMlo0I,
C_Din => CHTOLSRAML0Oi,
C_weN => CHTOLSRAMlL0l,
C_blK => "11",
C_wiDTH => CHTOLSRAMLoiL,
C_en => '1',
Sii_LOCk => '0',
BUsy => CHTOLSRAMl1OOl);
CHTOLSRAMlI0Ll: raM64x18
port map (A_doUT => CHTOLSRAMo1LI,
b_DOUt => open ,
A_addR_clk => Clk,
b_aDDR_cLK => CLK,
A_adDR_en => '1',
B_AddR_En => '1',
A_aDDR_laT => '1',
b_ADDr_LAT => '1',
A_addR_arsT_N => CHTOLSRAMil1,
B_addR_ArsT_N => CHTOLSRAMIl1,
a_ADdr_SRst_N => '1',
b_ADdr_SRst_N => '1',
A_DouT_Clk => '1',
b_DOUt_CLK => '1',
A_doUT_en => '1',
b_DOut_EN => '1',
A_dOUT_laT => '1',
b_DOut_LAt => '1',
A_dOUT_arST_n => CHTOLSRAMil1,
B_DouT_Arst_N => CHTOLSRAMIL1,
a_DOUt_SRSt_n => '1',
B_doUT_sRst_N => '1',
a_ADdr => CHTOLSRAMOL1i,
b_ADdr => CHTOLSRAMOl1i,
a_WidtH => CHTOLSRAMOoiL,
b_WidtH => CHTOLSRAMoOIl,
A_blK => CHTOLSRAMI111,
b_BLK => CHTOLSRAMoOOOl,
a_eN => '1',
b_EN => '1',
c_CLK => CLk,
C_AddR => CHTOLSRAMOO0i,
C_dIN => CHTOLSRAMO0oi,
C_weN => CHTOLSRAMOL0l,
C_bLK => "11",
c_WIdth => CHTOLSRAMoOIL,
C_en => '1',
Sii_LOck => '0',
busY => CHTOLSRAMi1oOL);
CHTOLSRAMIi0lL: RAm64X18
port map (a_DOut => CHTOLSRAMI0li,
B_doUT => open ,
A_adDR_clK => CLK,
b_Addr_CLk => clk,
a_aDDR_en => '1',
b_aDDr_eN => '1',
a_Addr_LAt => '1',
b_aDDr_lAT => '1',
A_adDR_arsT_n => CHTOLSRAMiL1,
B_adDR_arST_n => CHTOLSRAMIl1,
a_ADdr_SRSt_n => '1',
B_Addr_Srst_N => '1',
A_DouT_Clk => '1',
b_DOUt_CLK => '1',
A_dOUT_en => '1',
b_Dout_EN => '1',
a_DOUt_LAT => '1',
B_doUT_laT => '1',
a_Dout_ARst_N => CHTOLSRAMIL1,
b_DOUt_ARSt_n => CHTOLSRAMiL1,
A_doUT_srST_n => '1',
B_Dout_Srst_N => '1',
A_adDR => CHTOLSRAMio1I,
b_Addr => CHTOLSRAMIO1i,
A_wIDTh => CHTOLSRAMI1ll,
b_wIDTh => CHTOLSRAMI1lL,
a_BLk => CHTOLSRAMI111,
b_bLK => CHTOLSRAMOOool,
a_EN => '1',
b_EN => '1',
c_CLk => clk,
C_adDR => CHTOLSRAMi1iI,
c_DIn => CHTOLSRAMIIOi,
C_weN => CHTOLSRAMIO0l,
c_bLK => "11",
c_WidtH => CHTOLSRAMi1Ll,
C_en => '1',
SIi_lOCk => '0',
bUSY => CHTOLSRAMoOLOl);
CHTOLSRAMO00ll: rAM64x18
port map (A_Dout => CHTOLSRAMl0LI,
b_DOUt => open ,
A_Addr_Clk => cLK,
b_Addr_CLk => clK,
a_ADdr_EN => '1',
B_addR_En => '1',
a_aDDR_lAT => '1',
b_ADDr_lAT => '1',
A_Addr_Arst_N => CHTOLSRAMIl1,
b_aDDR_aRST_n => CHTOLSRAMil1,
a_aDDR_sRST_n => '1',
b_ADdr_SRSt_n => '1',
A_Dout_Clk => '1',
b_DOUt_CLK => '1',
A_douT_En => '1',
B_doUT_en => '1',
a_DOut_LAt => '1',
B_dOUT_laT => '1',
a_Dout_ARst_N => CHTOLSRAMIL1,
b_DOUt_ARSt_n => CHTOLSRAMil1,
A_doUT_srST_n => '1',
b_DOut_SRSt_n => '1',
a_aDDR => CHTOLSRAMlo1I,
B_AddR => CHTOLSRAMlO1I,
a_wIDTh => WIDth2,
B_wIDTh => WidtH2,
a_BLk => CHTOLSRAMI111,
B_blK => CHTOLSRAMoOOOl,
a_EN => '1',
B_eN => '1',
C_clK => cLK,
c_ADdr => CHTOLSRAML1ii,
c_DIN => CHTOLSRAMLIOi,
C_weN => CHTOLSRAMLO0l,
C_bLK => "11",
c_WIDth => wIDTh2,
c_EN => '1',
sII_locK => '0',
bUSY => CHTOLSRAMloLOL);
CHTOLSRAMl00Ll: raM64x18
port map (a_DOut => CHTOLSRAMO0li,
B_doUT => open ,
a_ADdr_CLk => cLK,
B_Addr_Clk => CLK,
A_adDR_en => '1',
b_ADdr_EN => '1',
A_addR_Lat => '1',
B_adDR_laT => '1',
a_Addr_ARst_N => CHTOLSRAMil1,
B_addR_arsT_N => CHTOLSRAMil1,
A_addR_srsT_N => '1',
b_ADdr_SRst_N => '1',
A_douT_Clk => '1',
b_DOUt_cLK => '1',
A_douT_En => '1',
b_DOUt_eN => '1',
A_douT_lat => '1',
b_DOut_LAt => '1',
a_DOUt_aRSt_n => CHTOLSRAMiL1,
B_dOUT_arST_n => CHTOLSRAMIl1,
a_DOut_SRst_N => '1',
b_dOUT_srST_n => '1',
a_ADdr => CHTOLSRAMOo1i,
b_Addr => CHTOLSRAMoo1I,
A_widTH => wiDTh1,
B_wIDTh => WIDth1,
a_bLK => CHTOLSRAMI111,
b_BLk => CHTOLSRAMoooOL,
A_en => '1',
B_en => '1',
c_cLK => CLk,
C_adDR => CHTOLSRAMO1iI,
c_DIn => CHTOLSRAMOIOi,
C_weN => CHTOLSRAMOo0l,
c_BLK => "11",
C_widTH => wiDTH1,
C_en => '1',
sii_Lock => '0',
busY => CHTOLSRAMIOLol);
CHTOLSRAMi00ll: rAM64x18
port map (a_Dout => CHTOLSRAMiiLI,
b_Dout => open ,
A_adDR_clk => CLk,
B_addR_Clk => cLK,
A_addR_en => '1',
b_ADDr_eN => '1',
A_adDR_laT => '1',
B_AddR_Lat => '1',
A_adDR_arsT_N => CHTOLSRAMIl1,
B_addR_ArsT_N => CHTOLSRAMIl1,
a_Addr_SRst_N => '1',
b_aDDr_sRST_n => '1',
A_DouT_Clk => '1',
B_douT_clk => '1',
a_DOut_EN => '1',
B_doUT_en => '1',
A_douT_Lat => '1',
b_Dout_LAt => '1',
a_DOUt_aRSt_n => CHTOLSRAMIL1,
b_dOUt_aRST_n => CHTOLSRAMiL1,
a_DOut_SRSt_n => '1',
B_doUT_srST_n => '1',
A_adDR => CHTOLSRAMi10I,
b_Addr => CHTOLSRAMi10I,
A_wiDTh => WidtH0,
B_WidTH => WIdth0,
a_BLk => CHTOLSRAMI111,
B_blK => CHTOLSRAMOOOol,
a_EN => '1',
B_en => '1',
C_clk => clK,
c_ADDr => CHTOLSRAMI0ii,
c_dIN => CHTOLSRAMILOi,
C_weN => CHTOLSRAMi1Il,
C_blK => "11",
c_wIDTh => WidTH0,
C_En => '1',
SII_loCK => '0',
buSY => CHTOLSRAMOLlol);
CHTOLSRAMLlloL <= CHTOLSRAMOLLol or CHTOLSRAMiOLOl
or CHTOLSRAMlolOL
or CHTOLSRAMOOLol
or CHTOLSRAMI1ooL
or CHTOLSRAML1Ool
or CHTOLSRAMo1oOL
or CHTOLSRAMI0ool
or CHTOLSRAMl0OOl
or CHTOLSRAMO0ooL
or CHTOLSRAMIIool
or CHTOLSRAMlIOOl
or CHTOLSRAMOiooL
or CHTOLSRAMiloOL
or CHTOLSRAMlLOOl
or CHTOLSRAMoloOL
or CHTOLSRAMLOooL
or CHTOLSRAMIoooL;
end architecture CHTOLSRAMo;
